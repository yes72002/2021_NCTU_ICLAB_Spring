`include "../00_TESTBED/pseudo_DRAM.sv"
`include "Usertype_PKG.sv"
`include "success.sv"
program automatic PATTERN(input clk, INF.PATTERN inf);
import usertype::*;

//================================================================
// parameters & integer
//================================================================
parameter DRAM_p_r = "../00_TESTBED/DRAM/dram.dat";
integer   wait_val_time, total_latency;
integer   lat;

//================================================================
// wire & registers 
//================================================================
logic [7:0] golden_DRAM[ ((65536+256*4)-1) : (65536+0) ];
// 10000(65536) ~ 103FC(66556)

Land_Info  golden_land_info;
Land       golden_land_id;
Crop_cat   golden_land_crop;
Crop_sta   golden_land_status;
Water_amnt golden_land_water;

logic      golden_complete;
Error_Msg  golden_err_msg;
logic [31:0] golden_deposit;
logic [31:0] golden_out_info;
logic [31:0] golden_out_deposit;

logic [7:0] golden_id;
// logic [3:0] golden_act;
Action      golden_act;
// logic [3:0] golden_crop;
Crop_cat golden_crop;
logic [15:0] golden_water;

//================================================================
// class random
//================================================================
class random_id;
        randc logic [7:0] ran_id;
        logic [7:0] ran_id_0  ;
		logic [7:0] out;
		// function new (int seed);
			// this.srandom(seed);
		// endfunction
        constraint range{ ran_id inside{[0:255]}; }
        // constraint range{ ran_id_0 inside{0}; }
		task set (logic [7:0] in);
			out = in;
		endtask
endclass

class random_act;
        rand Action ran_act;
        constraint range{ ran_act inside{Seed,Water,Reap,Steal}; }
endclass

class random_user_act_cnt;
        rand integer    ran_act_cnt;
        constraint range{ ran_act_cnt inside{[1:100]}; }
endclass

class random_crop;
        rand logic [3:0] ran_crop;
        constraint range{ ran_crop inside{Potato,Corn,Tomato,Wheat}; }
endclass

class random_water;
        rand logic [15:0] ran_water;
		rand logic [15:0] ran_water_0;
        rand logic [15:0] ran_water_1;
        rand logic [15:0] ran_water_2;
        rand logic [15:0] ran_water_3;
        rand logic [15:0] ran_water_4;
        rand logic [15:0] ran_water_5;
        constraint range{ ran_water inside{[0:1023]}; }
        constraint range_0{ ran_water_0 inside{[    0:12000]}; }
		constraint range_1{ ran_water_1 inside{[12001:24000]}; }
        constraint range_2{ ran_water_2 inside{[24001:36000]}; }
        constraint range_3{ ran_water_3 inside{[36001:48000]}; }
        constraint range_4{ ran_water_4 inside{[48001:60000]}; }
        constraint range_5{ ran_water_5 inside{[60001:65535]}; }
endclass


class random_passwd;
		rand logic [3:0]    ran_passwd;
		constraint range{ ran_passwd inside{[0:15]}; }
endclass


//================================================================
// initial
//================================================================
initial $readmemh(DRAM_p_r, golden_DRAM);
random_id            r_id      =  new();
random_act           r_act     =  new();
random_user_act_cnt  r_act_cnt =  new();
random_crop          r_crop    =  new();
random_water         r_water   =  new();
random_passwd        r_passwd  =  new();
initial begin
	inf.rst_n = 1;
	inf.id_valid = 0;
	inf.act_valid = 0;
	inf.cat_valid = 0;
	inf.amnt_valid = 0;
	inf.D = 'bx;
	
	golden_land_id = 0;
	golden_land_crop = 0;
	golden_land_status = 0;
	golden_land_water = 0;
	
	golden_err_msg = 0;
    golden_complete = 0;
	
	golden_id = 0;
	golden_act = 0;
	golden_crop = 0;
	golden_water = 0;
	
	golden_deposit  = 0;
	golden_out_info = 0;
	golden_out_deposit = 0;
	lat = 0;
	wait_val_time   = 0;
	total_latency   = 0;
	
	reset_signal_task;
	
	golden_deposit = {golden_DRAM[66556],golden_DRAM[66557],golden_DRAM[66558],golden_DRAM[66559]};
	
	// repeat(1) @(negedge clk);
	// give_check_deposit;
	// latency_task;
	// check_ans;
	
	give_id_0;
	// 1   - Seed
	// give_act_seed;
	give_act_seed_actual_0;	latency_task; check_ans;
	// 2   - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 3   - Water
	give_water_actual_0;	latency_task; check_ans;
	// 4   - Water
	give_water_actual_0;	latency_task; check_ans;
	// 5   - Reap
	give_act_reap;			latency_task; check_ans;
	// 6   - Reap
	give_act_reap;			latency_task; check_ans;
	// 7   - Steal
	give_act_steal;			latency_task; check_ans;
	// 8   - Steal
	give_act_steal;			latency_task; check_ans;
	// 9   - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 10  - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 11  - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 12  - Reap
	give_act_reap;			latency_task; check_ans;
	// 13  - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 14  - Water
	give_water_actual_0;	latency_task; check_ans;
	// 15  - Steal
	give_act_steal;			latency_task; check_ans;
	// 16  - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 17  - Steal
	give_act_steal;			latency_task; check_ans;
	// 18  - Water
	give_water_actual_0;	latency_task; check_ans;
	// 19  - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 20  - Reap
	give_act_reap;			latency_task; check_ans;
	// 21  - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 22  - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 23  - Steal
	give_act_steal;			latency_task; check_ans;
	// 24  - Reap
	give_act_reap;			latency_task; check_ans;
	// 25  - Water
	give_water_actual_0;	latency_task; check_ans;
	// 26  - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 27  - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 28  - Water
	give_water_actual_0;	latency_task; check_ans;
	// 29  - Water
	give_water_actual_0;	latency_task; check_ans;
	// 30  - Reap
	give_act_reap;			latency_task; check_ans;
	// 31  - Reap
	give_act_reap;			latency_task; check_ans;
	// 32  - Steal
	give_act_steal;			latency_task; check_ans;
	// 33  - Steal
	give_act_steal;			latency_task; check_ans;
	// 34  - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 35  - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 36  - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 37  - Reap
	give_act_reap;			latency_task; check_ans;
	// 38  - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 39  - Water
	give_water_actual_0;	latency_task; check_ans;
	// 40  - Steal
	give_act_steal;			latency_task; check_ans;
	// 41  - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 42  - Steal
	give_act_steal;			latency_task; check_ans;
	// 43  - Water
	give_water_actual_0;	latency_task; check_ans;
	// 44  - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 45  - Reap
	give_act_reap;			latency_task; check_ans;
	// 46  - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 47  - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 48  - Steal
	give_act_steal;			latency_task; check_ans;
	// 49  - Reap
	give_act_reap;			latency_task; check_ans;
	// 50  - Water
	give_water_actual_0;	latency_task; check_ans;
	// 51  - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 52  - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 53  - Water
	give_water_actual_0;	latency_task; check_ans;
	// 54  - Water
	give_water_actual_0;	latency_task; check_ans;
	// 55  - Reap
	give_act_reap;			latency_task; check_ans;
	// 56  - Reap
	give_act_reap;			latency_task; check_ans;
	// 57  - Steal
	give_act_steal;			latency_task; check_ans;
	// 58  - Steal
	give_act_steal;			latency_task; check_ans;
	// 59  - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 60  - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 61  - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 62  - Reap
	give_act_reap;			latency_task; check_ans;
	// 63  - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 64  - Water
	give_water_actual_0;	latency_task; check_ans;
	// 65  - Steal
	give_act_steal;			latency_task; check_ans;
	// 66  - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 67  - Steal
	give_act_steal;			latency_task; check_ans;
	// 68  - Water
	give_water_actual_0;	latency_task; check_ans;
	// 69  - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 70  - Reap
	give_act_reap;			latency_task; check_ans;
	// 71  - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 72  - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 73  - Steal
	give_act_steal;			latency_task; check_ans;
	// 74  - Reap
	give_act_reap;			latency_task; check_ans;
	// 75  - Water
	give_water_actual_0;	latency_task; check_ans;
	// 76  - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 77  - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 78  - Water
	give_water_actual_0;	latency_task; check_ans;
	// 79  - Water
	give_water_actual_0;	latency_task; check_ans;
	// 80  - Reap
	give_act_reap;			latency_task; check_ans;
	// 81  - Reap
	give_act_reap;			latency_task; check_ans;
	// 82  - Steal
	give_act_steal;			latency_task; check_ans;
	// 83  - Steal
	give_act_steal;			latency_task; check_ans;
	// 84  - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 85  - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 86  - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 87  - Reap
	give_act_reap;			latency_task; check_ans;
	// 88  - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 89  - Water
	give_water_actual_0;	latency_task; check_ans;
	// 90  - Steal
	give_act_steal;			latency_task; check_ans;
	// 91  - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 92  - Steal
	give_act_steal;			latency_task; check_ans;
	// 93  - Water
	give_water_actual_0;	latency_task; check_ans;
	// 94  - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 95  - Reap
	give_act_reap;			latency_task; check_ans;
	// 96  - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 97  - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 98  - Steal
	give_act_steal;			latency_task; check_ans;
	// 99  - Reap
	give_act_reap;			latency_task; check_ans;
	// 100 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 101 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 102 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 103 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 104 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 105 - Reap
	give_act_reap;			latency_task; check_ans;
	// 106 - Reap
	give_act_reap;			latency_task; check_ans;
	// 107 - Steal
	give_act_steal;			latency_task; check_ans;
	// 108 - Steal
	give_act_steal;			latency_task; check_ans;
	// 109 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 110 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 111 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 112 - Reap
	give_act_reap;			latency_task; check_ans;
	// 113 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 114 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 115 - Steal
	give_act_steal;			latency_task; check_ans;
	// 116 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 117 - Steal
	give_act_steal;			latency_task; check_ans;
	// 118 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 119 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 120 - Reap
	give_act_reap;			latency_task; check_ans;
	// 121 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 122 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 123 - Steal
	give_act_steal;			latency_task; check_ans;
	// 124 - Reap
	give_act_reap;			latency_task; check_ans;
	// 125 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 126 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 127 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 128 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 129 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 130 - Reap
	give_act_reap;			latency_task; check_ans;
	// 131 - Reap
	give_act_reap;			latency_task; check_ans;
	// 132 - Steal
	give_act_steal;			latency_task; check_ans;
	// 133 - Steal
	give_act_steal;			latency_task; check_ans;
	// 134 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 135 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 136 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 137 - Reap
	give_act_reap;			latency_task; check_ans;
	// 138 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 139 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 140 - Steal
	give_act_steal;			latency_task; check_ans;
	// 141 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 142 - Steal
	give_act_steal;			latency_task; check_ans;
	// 143 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 144 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 145 - Reap
	give_act_reap;			latency_task; check_ans;
	// 146 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 147 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 148 - Steal
	give_act_steal;			latency_task; check_ans;
	// 149 - Reap
	give_act_reap;			latency_task; check_ans;
	// 150 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 151 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 152 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 153 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 154 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 155 - Reap
	give_act_reap;			latency_task; check_ans;
	// 156 - Reap
	give_act_reap;			latency_task; check_ans;
	// 157 - Steal
	give_act_steal;			latency_task; check_ans;
	// 158 - Steal
	give_act_steal;			latency_task; check_ans;
	// 159 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 160 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 161 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 162 - Reap
	give_act_reap;			latency_task; check_ans;
	// 163 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 164 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 165 - Steal
	give_act_steal;			latency_task; check_ans;
	// 166 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 167 - Steal
	give_act_steal;			latency_task; check_ans;
	// 168 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 169 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 170 - Reap
	give_act_reap;			latency_task; check_ans;
	// 171 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 172 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 173 - Steal
	give_act_steal;			latency_task; check_ans;
	// 174 - Reap
	give_act_reap;			latency_task; check_ans;
	// 175 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 176 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 177 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 178 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 179 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 180 - Reap
	give_act_reap;			latency_task; check_ans;
	// 181 - Reap
	give_act_reap;			latency_task; check_ans;
	// 182 - Steal
	give_act_steal;			latency_task; check_ans;
	// 183 - Steal
	give_act_steal;			latency_task; check_ans;
	// 184 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 185 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 186 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 187 - Reap
	give_act_reap;			latency_task; check_ans;
	// 188 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 189 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 190 - Steal
	give_act_steal;			latency_task; check_ans;
	// 191 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 192 - Steal
	give_act_steal;			latency_task; check_ans;
	// 193 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 194 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 195 - Reap
	give_act_reap;			latency_task; check_ans;
	// 196 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 197 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 198 - Steal
	give_act_steal;			latency_task; check_ans;
	// 199 - Reap
	give_act_reap;			latency_task; check_ans;
	// 200 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 201 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 202 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 203 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 204 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 205 - Reap
	give_act_reap;			latency_task; check_ans;
	// 206 - Reap
	give_act_reap;			latency_task; check_ans;
	// 207 - Steal
	give_act_steal;			latency_task; check_ans;
	// 208 - Steal
	give_act_steal;			latency_task; check_ans;
	// 209 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 210 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 211 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 212 - Reap
	give_act_reap;			latency_task; check_ans;
	// 213 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 214 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 215 - Steal
	give_act_steal;			latency_task; check_ans;
	// 216 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 217 - Steal
	give_act_steal;			latency_task; check_ans;
	// 218 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 219 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 220 - Reap
	give_act_reap;			latency_task; check_ans;
	// 221 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 222 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 223 - Steal
	give_act_steal;			latency_task; check_ans;
	// 224 - Reap
	give_act_reap;			latency_task; check_ans;
	// 225 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 226 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 227 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 228 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 229 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 230 - Reap
	give_act_reap;			latency_task; check_ans;
	// 231 - Reap
	give_act_reap;			latency_task; check_ans;
	// 232 - Steal
	give_act_steal;			latency_task; check_ans;
	// 233 - Steal
	give_act_steal;			latency_task; check_ans;
	// 234 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 235 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 236 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 237 - Reap
	give_act_reap;			latency_task; check_ans;
	// 238 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 239 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 240 - Steal
	give_act_steal;			latency_task; check_ans;
	// 241 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 242 - Steal
	give_act_steal;			latency_task; check_ans;
	// 243 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 244 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 245 - Reap
	give_act_reap;			latency_task; check_ans;
	// 246 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	// 247 - Check_dep
	give_check_deposit;		latency_task; check_ans;
	// 248 - Steal
	give_act_steal;			latency_task; check_ans;
	// 249 - Reap
	give_act_reap;			latency_task; check_ans;
	// 250 - Water
	give_water_actual_0;	latency_task; check_ans;
	// 251 - Seed
	give_act_seed_actual_0;	latency_task; check_ans;
	
	// Spec 1 AMNT      20%
	// amnt1      100%  101
	// amnt2        0%    0
	// amnt3        0%    0
	// amnt4        0%    0
	// amnt5        0%    0
	// Spec 2 ID         0%
	// id[0]        0%    1
	// Spec 3 ACTION   100%
	// Spec 4 ERR_MSG   25%
	// Is_Empty     0%    0
	// Not_Empty    0%   50
	// Has_Grown    0%    0
	// Not_Grown  100%  100
	
	// 1 - Seed Water-amnt2
	give_act_seed_water_1; latency_task; check_ans;
	// 2  - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 3  - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 4  - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 5  - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 6  - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 7  - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 8  - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 9  - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 10 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 11 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 12 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 13 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 14 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 15 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 16 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 17 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 18 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 19 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 20 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 21 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 22 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 23 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 24 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 25 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 26 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 27 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 28 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 29 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 30 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 31 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 32 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 33 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 34 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 35 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 36 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 37 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 38 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 39 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 40 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 41 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 42 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 43 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 44 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 45 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 46 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 47 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 48 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 49 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	// 50 - Seed
	give_act_seed_water_1; latency_task; check_ans;
	
	// Spec 1 AMNT      20%
	// amnt1      100%  101
	// amnt2       50%   50
	// amnt3        0%    0
	// amnt4        0%    0
	// amnt5        0%    0
	// Spec 2 ID         0%
	// id[0]        0%    1
	// Spec 3 ACTION   100%
	// Spec 4 ERR_MSG   50%
	// Is_Empty     0%    0
	// Not_Empty  100%  100
	// Has_Grown    0%    0
	// Not_Grown  100%  100
	
	// 1   - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 2   - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 3   - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 4   - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 5   - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 6   - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 7   - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 8   - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 9   - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 10  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 11  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 12  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 13  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 14  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 15  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 16  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 17  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 18  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 19  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 20  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 21  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 22  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 23  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 24  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 25  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 26  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 27  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 28  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 29  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 30  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 31  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 32  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 33  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 34  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 35  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 36  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 37  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 38  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 39  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 40  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 41  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 42  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 43  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 44  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 45  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 46  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 47  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 48  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 49  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 50  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 51  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 52  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 53  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 54  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 55  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 56  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 57  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 58  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 59  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 60  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 61  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 62  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 63  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 64  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 65  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 66  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 67  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 68  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 69  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 70  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 71  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 72  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 73  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 74  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 75  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 76  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 77  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 78  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 79  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 80  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 81  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 82  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 83  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 84  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 85  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 86  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 87  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 88  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 89  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 90  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 91  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 92  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 93  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 94  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 95  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 96  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 97  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 98  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 99  - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 100 - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	// 101 - Water-amnt3 Has_Grown
	give_water_2; latency_task; check_ans;
	
	// Spec 1 AMNT      40%
	// amnt1      100%  101
	// amnt2       50%   50
	// amnt3      100%  101
	// amnt4        0%    0
	// amnt5        0%    0
	// Spec 2 ID         0%
	// id[0]        0%    1
	// Spec 3 ACTION   100%
	// Spec 4 ERR_MSG   75%
	// Is_Empty     0%    0
	// Not_Empty  100%  100
	// Has_Grown  100%  100
	// Not_Grown  100%  100

	// ID Water-amnt2 Is_Empty
	give_id_1  ; give_water_1; latency_task; check_ans;
	give_id_2  ; give_water_1; latency_task; check_ans;
	give_id_3  ; give_water_1; latency_task; check_ans;
	give_id_4  ; give_water_1; latency_task; check_ans;
	give_id_5  ; give_water_1; latency_task; check_ans;
	give_id_6  ; give_water_1; latency_task; check_ans;
	give_id_7  ; give_water_1; latency_task; check_ans;
	give_id_8  ; give_water_1; latency_task; check_ans;
	give_id_9  ; give_water_1; latency_task; check_ans;
	give_id_10 ; give_water_1; latency_task; check_ans;
	give_id_11 ; give_water_1; latency_task; check_ans;
	give_id_12 ; give_water_1; latency_task; check_ans;
	give_id_13 ; give_water_1; latency_task; check_ans;
	give_id_14 ; give_water_1; latency_task; check_ans;
	give_id_15 ; give_water_1; latency_task; check_ans;
	give_id_16 ; give_water_1; latency_task; check_ans;
	give_id_17 ; give_water_1; latency_task; check_ans;
	give_id_18 ; give_water_1; latency_task; check_ans;
	give_id_19 ; give_water_1; latency_task; check_ans;
	give_id_20 ; give_water_1; latency_task; check_ans;
	give_id_21 ; give_water_1; latency_task; check_ans;
	give_id_22 ; give_water_1; latency_task; check_ans;
	give_id_23 ; give_water_1; latency_task; check_ans;
	give_id_24 ; give_water_1; latency_task; check_ans;
	give_id_25 ; give_water_1; latency_task; check_ans;
	give_id_26 ; give_water_1; latency_task; check_ans;
	give_id_27 ; give_water_1; latency_task; check_ans;
	give_id_28 ; give_water_1; latency_task; check_ans;
	give_id_29 ; give_water_1; latency_task; check_ans;
	give_id_30 ; give_water_1; latency_task; check_ans;
	give_id_31 ; give_water_1; latency_task; check_ans;
	give_id_32 ; give_water_1; latency_task; check_ans;
	give_id_33 ; give_water_1; latency_task; check_ans;
	give_id_34 ; give_water_1; latency_task; check_ans;
	give_id_35 ; give_water_1; latency_task; check_ans;
	give_id_36 ; give_water_1; latency_task; check_ans;
	give_id_37 ; give_water_1; latency_task; check_ans;
	give_id_38 ; give_water_1; latency_task; check_ans;
	give_id_39 ; give_water_1; latency_task; check_ans;
	give_id_40 ; give_water_1; latency_task; check_ans;
	give_id_41 ; give_water_1; latency_task; check_ans;
	give_id_42 ; give_water_1; latency_task; check_ans;
	give_id_43 ; give_water_1; latency_task; check_ans;
	give_id_44 ; give_water_1; latency_task; check_ans;
	give_id_45 ; give_water_1; latency_task; check_ans;
	give_id_46 ; give_water_1; latency_task; check_ans;
	give_id_47 ; give_water_1; latency_task; check_ans;
	give_id_48 ; give_water_1; latency_task; check_ans;
	give_id_49 ; give_water_1; latency_task; check_ans;
	give_id_50 ; give_water_1; latency_task; check_ans;
	
	// Spec 1 AMNT      60%
	// amnt1      100%  101
	// amnt2      100%  100
	// amnt3      100%  101
	// amnt4        0%    0
	// amnt5        0%    0
	// Spec 2 ID         0%
	// id[0]        0%    1
	// Spec 3 ACTION   100%
	// Spec 4 ERR_MSG   75%
	// Is_Empty    50%   50
	// Not_Empty  100%  100
	// Has_Grown  100%  100
	// Not_Grown  100%  100
	
	// ID Water-amnt4 Is_Empty
	give_id_51 ; give_water_3; latency_task; check_ans;
	give_id_52 ; give_water_3; latency_task; check_ans;
	give_id_53 ; give_water_3; latency_task; check_ans;
	give_id_54 ; give_water_3; latency_task; check_ans;
	give_id_55 ; give_water_3; latency_task; check_ans;
	give_id_56 ; give_water_3; latency_task; check_ans;
	give_id_57 ; give_water_3; latency_task; check_ans;
	give_id_58 ; give_water_3; latency_task; check_ans;
	give_id_59 ; give_water_3; latency_task; check_ans;
	give_id_60 ; give_water_3; latency_task; check_ans;
	give_id_61 ; give_water_3; latency_task; check_ans;
	give_id_62 ; give_water_3; latency_task; check_ans;
	give_id_63 ; give_water_3; latency_task; check_ans;
	give_id_64 ; give_water_3; latency_task; check_ans;
	give_id_65 ; give_water_3; latency_task; check_ans;
	give_id_66 ; give_water_3; latency_task; check_ans;
	give_id_67 ; give_water_3; latency_task; check_ans;
	give_id_68 ; give_water_3; latency_task; check_ans;
	give_id_69 ; give_water_3; latency_task; check_ans;
	give_id_70 ; give_water_3; latency_task; check_ans;
	give_id_71 ; give_water_3; latency_task; check_ans;
	give_id_72 ; give_water_3; latency_task; check_ans;
	give_id_73 ; give_water_3; latency_task; check_ans;
	give_id_74 ; give_water_3; latency_task; check_ans;
	give_id_75 ; give_water_3; latency_task; check_ans;
	give_id_76 ; give_water_3; latency_task; check_ans;
	give_id_77 ; give_water_3; latency_task; check_ans;
	give_id_78 ; give_water_3; latency_task; check_ans;
	give_id_79 ; give_water_3; latency_task; check_ans;
	give_id_80 ; give_water_3; latency_task; check_ans;
	give_id_81 ; give_water_3; latency_task; check_ans;
	give_id_82 ; give_water_3; latency_task; check_ans;
	give_id_83 ; give_water_3; latency_task; check_ans;
	give_id_84 ; give_water_3; latency_task; check_ans;
	give_id_85 ; give_water_3; latency_task; check_ans;
	give_id_86 ; give_water_3; latency_task; check_ans;
	give_id_87 ; give_water_3; latency_task; check_ans;
	give_id_88 ; give_water_3; latency_task; check_ans;
	give_id_89 ; give_water_3; latency_task; check_ans;
	give_id_90 ; give_water_3; latency_task; check_ans;
	give_id_91 ; give_water_3; latency_task; check_ans;
	give_id_92 ; give_water_3; latency_task; check_ans;
	give_id_93 ; give_water_3; latency_task; check_ans;
	give_id_94 ; give_water_3; latency_task; check_ans;
	give_id_95 ; give_water_3; latency_task; check_ans;
	give_id_96 ; give_water_3; latency_task; check_ans;
	give_id_97 ; give_water_3; latency_task; check_ans;
	give_id_98 ; give_water_3; latency_task; check_ans;
	give_id_99 ; give_water_3; latency_task; check_ans;
	give_id_100; give_water_3; latency_task; check_ans;
	give_id_101; give_water_3; latency_task; check_ans;
	give_id_102; give_water_3; latency_task; check_ans;
	give_id_103; give_water_3; latency_task; check_ans;
	give_id_104; give_water_3; latency_task; check_ans;
	give_id_105; give_water_3; latency_task; check_ans;
	give_id_106; give_water_3; latency_task; check_ans;
	give_id_107; give_water_3; latency_task; check_ans;
	give_id_108; give_water_3; latency_task; check_ans;
	give_id_109; give_water_3; latency_task; check_ans;
	give_id_110; give_water_3; latency_task; check_ans;
	give_id_111; give_water_3; latency_task; check_ans;
	give_id_112; give_water_3; latency_task; check_ans;
	give_id_113; give_water_3; latency_task; check_ans;
	give_id_114; give_water_3; latency_task; check_ans;
	give_id_115; give_water_3; latency_task; check_ans;
	give_id_116; give_water_3; latency_task; check_ans;
	give_id_117; give_water_3; latency_task; check_ans;
	give_id_118; give_water_3; latency_task; check_ans;
	give_id_119; give_water_3; latency_task; check_ans;
	give_id_120; give_water_3; latency_task; check_ans;
	give_id_121; give_water_3; latency_task; check_ans;
	give_id_122; give_water_3; latency_task; check_ans;
	give_id_123; give_water_3; latency_task; check_ans;
	give_id_124; give_water_3; latency_task; check_ans;
	give_id_125; give_water_3; latency_task; check_ans;
	give_id_126; give_water_3; latency_task; check_ans;
	give_id_127; give_water_3; latency_task; check_ans;
	give_id_128; give_water_3; latency_task; check_ans;
	give_id_129; give_water_3; latency_task; check_ans;
	give_id_130; give_water_3; latency_task; check_ans;
	give_id_131; give_water_3; latency_task; check_ans;
	give_id_132; give_water_3; latency_task; check_ans;
	give_id_133; give_water_3; latency_task; check_ans;
	give_id_134; give_water_3; latency_task; check_ans;
	give_id_135; give_water_3; latency_task; check_ans;
	give_id_136; give_water_3; latency_task; check_ans;
	give_id_137; give_water_3; latency_task; check_ans;
	give_id_138; give_water_3; latency_task; check_ans;
	give_id_139; give_water_3; latency_task; check_ans;
	give_id_140; give_water_3; latency_task; check_ans;
	give_id_141; give_water_3; latency_task; check_ans;
	give_id_142; give_water_3; latency_task; check_ans;
	give_id_143; give_water_3; latency_task; check_ans;
	give_id_144; give_water_3; latency_task; check_ans;
	give_id_145; give_water_3; latency_task; check_ans;
	give_id_146; give_water_3; latency_task; check_ans;
	give_id_147; give_water_3; latency_task; check_ans;
	give_id_148; give_water_3; latency_task; check_ans;
	give_id_149; give_water_3; latency_task; check_ans;
	give_id_150; give_water_3; latency_task; check_ans;
	
	// Spec 1 AMNT      80%
	// amnt1      100%  101
	// amnt2      100%  100
	// amnt3      100%  101
	// amnt4      100%  100
	// amnt5        0%    0
	// Spec 2 ID         0%
	// id[0]        0%    1
	// Spec 3 ACTION   100%
	// Spec 4 ERR_MSG  100%
	// Is_Empty   100%  150
	// Not_Empty  100%  100
	// Has_Grown  100%  100
	// Not_Grown  100%  100
	
	// ID Water-amnt5 Is_Empty
	give_id_151; give_water_4; latency_task; check_ans;
	give_id_152; give_water_4; latency_task; check_ans;
	give_id_153; give_water_4; latency_task; check_ans;
	give_id_154; give_water_4; latency_task; check_ans;
	give_id_155; give_water_4; latency_task; check_ans;
	give_id_156; give_water_4; latency_task; check_ans;
	give_id_157; give_water_4; latency_task; check_ans;
	give_id_158; give_water_4; latency_task; check_ans;
	give_id_159; give_water_4; latency_task; check_ans;
	give_id_160; give_water_4; latency_task; check_ans;
	give_id_161; give_water_4; latency_task; check_ans;
	give_id_162; give_water_4; latency_task; check_ans;
	give_id_163; give_water_4; latency_task; check_ans;
	give_id_164; give_water_4; latency_task; check_ans;
	give_id_165; give_water_4; latency_task; check_ans;
	give_id_166; give_water_4; latency_task; check_ans;
	give_id_167; give_water_4; latency_task; check_ans;
	give_id_168; give_water_4; latency_task; check_ans;
	give_id_169; give_water_4; latency_task; check_ans;
	give_id_170; give_water_4; latency_task; check_ans;
	give_id_171; give_water_4; latency_task; check_ans;
	give_id_172; give_water_4; latency_task; check_ans;
	give_id_173; give_water_4; latency_task; check_ans;
	give_id_174; give_water_4; latency_task; check_ans;
	give_id_175; give_water_4; latency_task; check_ans;
	give_id_176; give_water_4; latency_task; check_ans;
	give_id_177; give_water_4; latency_task; check_ans;
	give_id_178; give_water_4; latency_task; check_ans;
	give_id_179; give_water_4; latency_task; check_ans;
	give_id_180; give_water_4; latency_task; check_ans;
	give_id_181; give_water_4; latency_task; check_ans;
	give_id_182; give_water_4; latency_task; check_ans;
	give_id_183; give_water_4; latency_task; check_ans;
	give_id_184; give_water_4; latency_task; check_ans;
	give_id_185; give_water_4; latency_task; check_ans;
	give_id_186; give_water_4; latency_task; check_ans;
	give_id_187; give_water_4; latency_task; check_ans;
	give_id_188; give_water_4; latency_task; check_ans;
	give_id_189; give_water_4; latency_task; check_ans;
	give_id_190; give_water_4; latency_task; check_ans;
	give_id_191; give_water_4; latency_task; check_ans;
	give_id_192; give_water_4; latency_task; check_ans;
	give_id_193; give_water_4; latency_task; check_ans;
	give_id_194; give_water_4; latency_task; check_ans;
	give_id_195; give_water_4; latency_task; check_ans;
	give_id_196; give_water_4; latency_task; check_ans;
	give_id_197; give_water_4; latency_task; check_ans;
	give_id_198; give_water_4; latency_task; check_ans;
	give_id_199; give_water_4; latency_task; check_ans;
	give_id_200; give_water_4; latency_task; check_ans;
	give_id_201; give_water_4; latency_task; check_ans;
	give_id_202; give_water_4; latency_task; check_ans;
	give_id_203; give_water_4; latency_task; check_ans;
	give_id_204; give_water_4; latency_task; check_ans;
	give_id_205; give_water_4; latency_task; check_ans;
	give_id_206; give_water_4; latency_task; check_ans;
	give_id_207; give_water_4; latency_task; check_ans;
	give_id_208; give_water_4; latency_task; check_ans;
	give_id_209; give_water_4; latency_task; check_ans;
	give_id_210; give_water_4; latency_task; check_ans;
	give_id_211; give_water_4; latency_task; check_ans;
	give_id_212; give_water_4; latency_task; check_ans;
	give_id_213; give_water_4; latency_task; check_ans;
	give_id_214; give_water_4; latency_task; check_ans;
	give_id_215; give_water_4; latency_task; check_ans;
	give_id_216; give_water_4; latency_task; check_ans;
	give_id_217; give_water_4; latency_task; check_ans;
	give_id_218; give_water_4; latency_task; check_ans;
	give_id_219; give_water_4; latency_task; check_ans;
	give_id_220; give_water_4; latency_task; check_ans;
	give_id_221; give_water_4; latency_task; check_ans;
	give_id_222; give_water_4; latency_task; check_ans;
	give_id_223; give_water_4; latency_task; check_ans;
	give_id_224; give_water_4; latency_task; check_ans;
	give_id_225; give_water_4; latency_task; check_ans;
	give_id_226; give_water_4; latency_task; check_ans;
	give_id_227; give_water_4; latency_task; check_ans;
	give_id_228; give_water_4; latency_task; check_ans;
	give_id_229; give_water_4; latency_task; check_ans;
	give_id_230; give_water_4; latency_task; check_ans;
	give_id_231; give_water_4; latency_task; check_ans;
	give_id_232; give_water_4; latency_task; check_ans;
	give_id_233; give_water_4; latency_task; check_ans;
	give_id_234; give_water_4; latency_task; check_ans;
	give_id_235; give_water_4; latency_task; check_ans;
	give_id_236; give_water_4; latency_task; check_ans;
	give_id_237; give_water_4; latency_task; check_ans;
	give_id_238; give_water_4; latency_task; check_ans;
	give_id_239; give_water_4; latency_task; check_ans;
	give_id_240; give_water_4; latency_task; check_ans;
	give_id_241; give_water_4; latency_task; check_ans;
	give_id_242; give_water_4; latency_task; check_ans;
	give_id_243; give_water_4; latency_task; check_ans;
	give_id_244; give_water_4; latency_task; check_ans;
	give_id_245; give_water_4; latency_task; check_ans;
	give_id_246; give_water_4; latency_task; check_ans;
	give_id_247; give_water_4; latency_task; check_ans;
	give_id_248; give_water_4; latency_task; check_ans;
	give_id_249; give_water_4; latency_task; check_ans;
	give_id_250; give_water_4; latency_task; check_ans;
	give_id_251; give_water_4; latency_task; check_ans;
	give_id_252; give_water_4; latency_task; check_ans;
	give_id_253; give_water_4; latency_task; check_ans;
	give_id_254; give_water_4; latency_task; check_ans;

	// Spec 1 AMNT     100%
	// amnt1      100%  101
	// amnt2      100%  100
	// amnt3      100%  101
	// amnt4      100%  100
	// amnt5      100%  104
	// Spec 2 ID         0%
	// id[0]~id[254]0%    1
	// Spec 3 ACTION   100%
	// Spec 4 ERR_MSG  100%
	// Is_Empty   100%  254
	// Not_Empty  100%  100
	// Has_Grown  100%  100
	// Not_Grown  100%  100
	
	// give_id_0; give_water_4; latency_task; check_ans; //195620
	// give_id_0; give_act_reap; latency_task; check_ans; //195590
	// give_id_0; give_act_steal; latency_task; check_ans; //195590
	// give_id_0; give_check_deposit; latency_task; check_ans; //195590
	// ID 2
	give_id_0  ; give_act_reap; latency_task; check_ans;
	give_id_1  ; give_act_reap; latency_task; check_ans;
	give_id_2  ; give_act_reap; latency_task; check_ans;
	give_id_3  ; give_act_reap; latency_task; check_ans;
	give_id_4  ; give_act_reap; latency_task; check_ans;
	give_id_5  ; give_act_reap; latency_task; check_ans;
	give_id_6  ; give_act_reap; latency_task; check_ans;
	give_id_7  ; give_act_reap; latency_task; check_ans;
	give_id_8  ; give_act_reap; latency_task; check_ans;
	give_id_9  ; give_act_reap; latency_task; check_ans;
	give_id_10 ; give_act_reap; latency_task; check_ans;
	give_id_11 ; give_act_reap; latency_task; check_ans;
	give_id_12 ; give_act_reap; latency_task; check_ans;
	give_id_13 ; give_act_reap; latency_task; check_ans;
	give_id_14 ; give_act_reap; latency_task; check_ans;
	give_id_15 ; give_act_reap; latency_task; check_ans;
	give_id_16 ; give_act_reap; latency_task; check_ans;
	give_id_17 ; give_act_reap; latency_task; check_ans;
	give_id_18 ; give_act_reap; latency_task; check_ans;
	give_id_19 ; give_act_reap; latency_task; check_ans;
	give_id_20 ; give_act_reap; latency_task; check_ans;
	give_id_21 ; give_act_reap; latency_task; check_ans;
	give_id_22 ; give_act_reap; latency_task; check_ans;
	give_id_23 ; give_act_reap; latency_task; check_ans;
	give_id_24 ; give_act_reap; latency_task; check_ans;
	give_id_25 ; give_act_reap; latency_task; check_ans;
	give_id_26 ; give_act_reap; latency_task; check_ans;
	give_id_27 ; give_act_reap; latency_task; check_ans;
	give_id_28 ; give_act_reap; latency_task; check_ans;
	give_id_29 ; give_act_reap; latency_task; check_ans;
	give_id_30 ; give_act_reap; latency_task; check_ans;
	give_id_31 ; give_act_reap; latency_task; check_ans;
	give_id_32 ; give_act_reap; latency_task; check_ans;
	give_id_33 ; give_act_reap; latency_task; check_ans;
	give_id_34 ; give_act_reap; latency_task; check_ans;
	give_id_35 ; give_act_reap; latency_task; check_ans;
	give_id_36 ; give_act_reap; latency_task; check_ans;
	give_id_37 ; give_act_reap; latency_task; check_ans;
	give_id_38 ; give_act_reap; latency_task; check_ans;
	give_id_39 ; give_act_reap; latency_task; check_ans;
	give_id_40 ; give_act_reap; latency_task; check_ans;
	give_id_41 ; give_act_reap; latency_task; check_ans;
	give_id_42 ; give_act_reap; latency_task; check_ans;
	give_id_43 ; give_act_reap; latency_task; check_ans;
	give_id_44 ; give_act_reap; latency_task; check_ans;
	give_id_45 ; give_act_reap; latency_task; check_ans;
	give_id_46 ; give_act_reap; latency_task; check_ans;
	give_id_47 ; give_act_reap; latency_task; check_ans;
	give_id_48 ; give_act_reap; latency_task; check_ans;
	give_id_49 ; give_act_reap; latency_task; check_ans;
	give_id_50 ; give_act_reap; latency_task; check_ans;
	give_id_51 ; give_act_reap; latency_task; check_ans;
	give_id_52 ; give_act_reap; latency_task; check_ans;
	give_id_53 ; give_act_reap; latency_task; check_ans;
	give_id_54 ; give_act_reap; latency_task; check_ans;
	give_id_55 ; give_act_reap; latency_task; check_ans;
	give_id_56 ; give_act_reap; latency_task; check_ans;
	give_id_57 ; give_act_reap; latency_task; check_ans;
	give_id_58 ; give_act_reap; latency_task; check_ans;
	give_id_59 ; give_act_reap; latency_task; check_ans;
	give_id_60 ; give_act_reap; latency_task; check_ans;
	give_id_61 ; give_act_reap; latency_task; check_ans;
	give_id_62 ; give_act_reap; latency_task; check_ans;
	give_id_63 ; give_act_reap; latency_task; check_ans;
	give_id_64 ; give_act_reap; latency_task; check_ans;
	give_id_65 ; give_act_reap; latency_task; check_ans;
	give_id_66 ; give_act_reap; latency_task; check_ans;
	give_id_67 ; give_act_reap; latency_task; check_ans;
	give_id_68 ; give_act_reap; latency_task; check_ans;
	give_id_69 ; give_act_reap; latency_task; check_ans;
	give_id_70 ; give_act_reap; latency_task; check_ans;
	give_id_71 ; give_act_reap; latency_task; check_ans;
	give_id_72 ; give_act_reap; latency_task; check_ans;
	give_id_73 ; give_act_reap; latency_task; check_ans;
	give_id_74 ; give_act_reap; latency_task; check_ans;
	give_id_75 ; give_act_reap; latency_task; check_ans;
	give_id_76 ; give_act_reap; latency_task; check_ans;
	give_id_77 ; give_act_reap; latency_task; check_ans;
	give_id_78 ; give_act_reap; latency_task; check_ans;
	give_id_79 ; give_act_reap; latency_task; check_ans;
	give_id_80 ; give_act_reap; latency_task; check_ans;
	give_id_81 ; give_act_reap; latency_task; check_ans;
	give_id_82 ; give_act_reap; latency_task; check_ans;
	give_id_83 ; give_act_reap; latency_task; check_ans;
	give_id_84 ; give_act_reap; latency_task; check_ans;
	give_id_85 ; give_act_reap; latency_task; check_ans;
	give_id_86 ; give_act_reap; latency_task; check_ans;
	give_id_87 ; give_act_reap; latency_task; check_ans;
	give_id_88 ; give_act_reap; latency_task; check_ans;
	give_id_89 ; give_act_reap; latency_task; check_ans;
	give_id_90 ; give_act_reap; latency_task; check_ans;
	give_id_91 ; give_act_reap; latency_task; check_ans;
	give_id_92 ; give_act_reap; latency_task; check_ans;
	give_id_93 ; give_act_reap; latency_task; check_ans;
	give_id_94 ; give_act_reap; latency_task; check_ans;
	give_id_95 ; give_act_reap; latency_task; check_ans;
	give_id_96 ; give_act_reap; latency_task; check_ans;
	give_id_97 ; give_act_reap; latency_task; check_ans;
	give_id_98 ; give_act_reap; latency_task; check_ans;
	give_id_99 ; give_act_reap; latency_task; check_ans;
	give_id_100; give_act_reap; latency_task; check_ans;
	give_id_101; give_act_reap; latency_task; check_ans;
	give_id_102; give_act_reap; latency_task; check_ans;
	give_id_103; give_act_reap; latency_task; check_ans;
	give_id_104; give_act_reap; latency_task; check_ans;
	give_id_105; give_act_reap; latency_task; check_ans;
	give_id_106; give_act_reap; latency_task; check_ans;
	give_id_107; give_act_reap; latency_task; check_ans;
	give_id_108; give_act_reap; latency_task; check_ans;
	give_id_109; give_act_reap; latency_task; check_ans;
	give_id_110; give_act_reap; latency_task; check_ans;
	give_id_111; give_act_reap; latency_task; check_ans;
	give_id_112; give_act_reap; latency_task; check_ans;
	give_id_113; give_act_reap; latency_task; check_ans;
	give_id_114; give_act_reap; latency_task; check_ans;
	give_id_115; give_act_reap; latency_task; check_ans;
	give_id_116; give_act_reap; latency_task; check_ans;
	give_id_117; give_act_reap; latency_task; check_ans;
	give_id_118; give_act_reap; latency_task; check_ans;
	give_id_119; give_act_reap; latency_task; check_ans;
	give_id_120; give_act_reap; latency_task; check_ans;
	give_id_121; give_act_reap; latency_task; check_ans;
	give_id_122; give_act_reap; latency_task; check_ans;
	give_id_123; give_act_reap; latency_task; check_ans;
	give_id_124; give_act_reap; latency_task; check_ans;
	give_id_125; give_act_reap; latency_task; check_ans;
	give_id_126; give_act_reap; latency_task; check_ans;
	give_id_127; give_act_reap; latency_task; check_ans;
	give_id_128; give_act_reap; latency_task; check_ans;
	give_id_129; give_act_reap; latency_task; check_ans;
	give_id_130; give_act_reap; latency_task; check_ans;
	give_id_131; give_act_reap; latency_task; check_ans;
	give_id_132; give_act_reap; latency_task; check_ans;
	give_id_133; give_act_reap; latency_task; check_ans;
	give_id_134; give_act_reap; latency_task; check_ans;
	give_id_135; give_act_reap; latency_task; check_ans;
	give_id_136; give_act_reap; latency_task; check_ans;
	give_id_137; give_act_reap; latency_task; check_ans;
	give_id_138; give_act_reap; latency_task; check_ans;
	give_id_139; give_act_reap; latency_task; check_ans;
	give_id_140; give_act_reap; latency_task; check_ans;
	give_id_141; give_act_reap; latency_task; check_ans;
	give_id_142; give_act_reap; latency_task; check_ans;
	give_id_143; give_act_reap; latency_task; check_ans;
	give_id_144; give_act_reap; latency_task; check_ans;
	give_id_145; give_act_reap; latency_task; check_ans;
	give_id_146; give_act_reap; latency_task; check_ans;
	give_id_147; give_act_reap; latency_task; check_ans;
	give_id_148; give_act_reap; latency_task; check_ans;
	give_id_149; give_act_reap; latency_task; check_ans;
	give_id_150; give_act_reap; latency_task; check_ans;
	give_id_151; give_act_reap; latency_task; check_ans;
	give_id_152; give_act_reap; latency_task; check_ans;
	give_id_153; give_act_reap; latency_task; check_ans;
	give_id_154; give_act_reap; latency_task; check_ans;
	give_id_155; give_act_reap; latency_task; check_ans;
	give_id_156; give_act_reap; latency_task; check_ans;
	give_id_157; give_act_reap; latency_task; check_ans;
	give_id_158; give_act_reap; latency_task; check_ans;
	give_id_159; give_act_reap; latency_task; check_ans;
	give_id_160; give_act_reap; latency_task; check_ans;
	give_id_161; give_act_reap; latency_task; check_ans;
	give_id_162; give_act_reap; latency_task; check_ans;
	give_id_163; give_act_reap; latency_task; check_ans;
	give_id_164; give_act_reap; latency_task; check_ans;
	give_id_165; give_act_reap; latency_task; check_ans;
	give_id_166; give_act_reap; latency_task; check_ans;
	give_id_167; give_act_reap; latency_task; check_ans;
	give_id_168; give_act_reap; latency_task; check_ans;
	give_id_169; give_act_reap; latency_task; check_ans;
	give_id_170; give_act_reap; latency_task; check_ans;
	give_id_171; give_act_reap; latency_task; check_ans;
	give_id_172; give_act_reap; latency_task; check_ans;
	give_id_173; give_act_reap; latency_task; check_ans;
	give_id_174; give_act_reap; latency_task; check_ans;
	give_id_175; give_act_reap; latency_task; check_ans;
	give_id_176; give_act_reap; latency_task; check_ans;
	give_id_177; give_act_reap; latency_task; check_ans;
	give_id_178; give_act_reap; latency_task; check_ans;
	give_id_179; give_act_reap; latency_task; check_ans;
	give_id_180; give_act_reap; latency_task; check_ans;
	give_id_181; give_act_reap; latency_task; check_ans;
	give_id_182; give_act_reap; latency_task; check_ans;
	give_id_183; give_act_reap; latency_task; check_ans;
	give_id_184; give_act_reap; latency_task; check_ans;
	give_id_185; give_act_reap; latency_task; check_ans;
	give_id_186; give_act_reap; latency_task; check_ans;
	give_id_187; give_act_reap; latency_task; check_ans;
	give_id_188; give_act_reap; latency_task; check_ans;
	give_id_189; give_act_reap; latency_task; check_ans;
	give_id_190; give_act_reap; latency_task; check_ans;
	give_id_191; give_act_reap; latency_task; check_ans;
	give_id_192; give_act_reap; latency_task; check_ans;
	give_id_193; give_act_reap; latency_task; check_ans;
	give_id_194; give_act_reap; latency_task; check_ans;
	give_id_195; give_act_reap; latency_task; check_ans;
	give_id_196; give_act_reap; latency_task; check_ans;
	give_id_197; give_act_reap; latency_task; check_ans;
	give_id_198; give_act_reap; latency_task; check_ans;
	give_id_199; give_act_reap; latency_task; check_ans;
	give_id_200; give_act_reap; latency_task; check_ans;
	give_id_201; give_act_reap; latency_task; check_ans;
	give_id_202; give_act_reap; latency_task; check_ans;
	give_id_203; give_act_reap; latency_task; check_ans;
	give_id_204; give_act_reap; latency_task; check_ans;
	give_id_205; give_act_reap; latency_task; check_ans;
	give_id_206; give_act_reap; latency_task; check_ans;
	give_id_207; give_act_reap; latency_task; check_ans;
	give_id_208; give_act_reap; latency_task; check_ans;
	give_id_209; give_act_reap; latency_task; check_ans;
	give_id_210; give_act_reap; latency_task; check_ans;
	give_id_211; give_act_reap; latency_task; check_ans;
	give_id_212; give_act_reap; latency_task; check_ans;
	give_id_213; give_act_reap; latency_task; check_ans;
	give_id_214; give_act_reap; latency_task; check_ans;
	give_id_215; give_act_reap; latency_task; check_ans;
	give_id_216; give_act_reap; latency_task; check_ans;
	give_id_217; give_act_reap; latency_task; check_ans;
	give_id_218; give_act_reap; latency_task; check_ans;
	give_id_219; give_act_reap; latency_task; check_ans;
	give_id_220; give_act_reap; latency_task; check_ans;
	give_id_221; give_act_reap; latency_task; check_ans;
	give_id_222; give_act_reap; latency_task; check_ans;
	give_id_223; give_act_reap; latency_task; check_ans;
	give_id_224; give_act_reap; latency_task; check_ans;
	give_id_225; give_act_reap; latency_task; check_ans;
	give_id_226; give_act_reap; latency_task; check_ans;
	give_id_227; give_act_reap; latency_task; check_ans;
	give_id_228; give_act_reap; latency_task; check_ans;
	give_id_229; give_act_reap; latency_task; check_ans;
	give_id_230; give_act_reap; latency_task; check_ans;
	give_id_231; give_act_reap; latency_task; check_ans;
	give_id_232; give_act_reap; latency_task; check_ans;
	give_id_233; give_act_reap; latency_task; check_ans;
	give_id_234; give_act_reap; latency_task; check_ans;
	give_id_235; give_act_reap; latency_task; check_ans;
	give_id_236; give_act_reap; latency_task; check_ans;
	give_id_237; give_act_reap; latency_task; check_ans;
	give_id_238; give_act_reap; latency_task; check_ans;
	give_id_239; give_act_reap; latency_task; check_ans;
	give_id_240; give_act_reap; latency_task; check_ans;
	give_id_241; give_act_reap; latency_task; check_ans;
	give_id_242; give_act_reap; latency_task; check_ans;
	give_id_243; give_act_reap; latency_task; check_ans;
	give_id_244; give_act_reap; latency_task; check_ans;
	give_id_245; give_act_reap; latency_task; check_ans;
	give_id_246; give_act_reap; latency_task; check_ans;
	give_id_247; give_act_reap; latency_task; check_ans;
	give_id_248; give_act_reap; latency_task; check_ans;
	give_id_249; give_act_reap; latency_task; check_ans;
	give_id_250; give_act_reap; latency_task; check_ans;
	give_id_251; give_act_reap; latency_task; check_ans;
	give_id_252; give_act_reap; latency_task; check_ans;
	give_id_253; give_act_reap; latency_task; check_ans;
	give_id_254; give_act_reap; latency_task; check_ans;
	// ID 3
	give_id_0  ; give_act_reap; latency_task; check_ans;
	give_id_1  ; give_act_reap; latency_task; check_ans;
	give_id_2  ; give_act_reap; latency_task; check_ans;
	give_id_3  ; give_act_reap; latency_task; check_ans;
	give_id_4  ; give_act_reap; latency_task; check_ans;
	give_id_5  ; give_act_reap; latency_task; check_ans;
	give_id_6  ; give_act_reap; latency_task; check_ans;
	give_id_7  ; give_act_reap; latency_task; check_ans;
	give_id_8  ; give_act_reap; latency_task; check_ans;
	give_id_9  ; give_act_reap; latency_task; check_ans;
	give_id_10 ; give_act_reap; latency_task; check_ans;
	give_id_11 ; give_act_reap; latency_task; check_ans;
	give_id_12 ; give_act_reap; latency_task; check_ans;
	give_id_13 ; give_act_reap; latency_task; check_ans;
	give_id_14 ; give_act_reap; latency_task; check_ans;
	give_id_15 ; give_act_reap; latency_task; check_ans;
	give_id_16 ; give_act_reap; latency_task; check_ans;
	give_id_17 ; give_act_reap; latency_task; check_ans;
	give_id_18 ; give_act_reap; latency_task; check_ans;
	give_id_19 ; give_act_reap; latency_task; check_ans;
	give_id_20 ; give_act_reap; latency_task; check_ans;
	give_id_21 ; give_act_reap; latency_task; check_ans;
	give_id_22 ; give_act_reap; latency_task; check_ans;
	give_id_23 ; give_act_reap; latency_task; check_ans;
	give_id_24 ; give_act_reap; latency_task; check_ans;
	give_id_25 ; give_act_reap; latency_task; check_ans;
	give_id_26 ; give_act_reap; latency_task; check_ans;
	give_id_27 ; give_act_reap; latency_task; check_ans;
	give_id_28 ; give_act_reap; latency_task; check_ans;
	give_id_29 ; give_act_reap; latency_task; check_ans;
	give_id_30 ; give_act_reap; latency_task; check_ans;
	give_id_31 ; give_act_reap; latency_task; check_ans;
	give_id_32 ; give_act_reap; latency_task; check_ans;
	give_id_33 ; give_act_reap; latency_task; check_ans;
	give_id_34 ; give_act_reap; latency_task; check_ans;
	give_id_35 ; give_act_reap; latency_task; check_ans;
	give_id_36 ; give_act_reap; latency_task; check_ans;
	give_id_37 ; give_act_reap; latency_task; check_ans;
	give_id_38 ; give_act_reap; latency_task; check_ans;
	give_id_39 ; give_act_reap; latency_task; check_ans;
	give_id_40 ; give_act_reap; latency_task; check_ans;
	give_id_41 ; give_act_reap; latency_task; check_ans;
	give_id_42 ; give_act_reap; latency_task; check_ans;
	give_id_43 ; give_act_reap; latency_task; check_ans;
	give_id_44 ; give_act_reap; latency_task; check_ans;
	give_id_45 ; give_act_reap; latency_task; check_ans;
	give_id_46 ; give_act_reap; latency_task; check_ans;
	give_id_47 ; give_act_reap; latency_task; check_ans;
	give_id_48 ; give_act_reap; latency_task; check_ans;
	give_id_49 ; give_act_reap; latency_task; check_ans;
	give_id_50 ; give_act_reap; latency_task; check_ans;
	give_id_51 ; give_act_reap; latency_task; check_ans;
	give_id_52 ; give_act_reap; latency_task; check_ans;
	give_id_53 ; give_act_reap; latency_task; check_ans;
	give_id_54 ; give_act_reap; latency_task; check_ans;
	give_id_55 ; give_act_reap; latency_task; check_ans;
	give_id_56 ; give_act_reap; latency_task; check_ans;
	give_id_57 ; give_act_reap; latency_task; check_ans;
	give_id_58 ; give_act_reap; latency_task; check_ans;
	give_id_59 ; give_act_reap; latency_task; check_ans;
	give_id_60 ; give_act_reap; latency_task; check_ans;
	give_id_61 ; give_act_reap; latency_task; check_ans;
	give_id_62 ; give_act_reap; latency_task; check_ans;
	give_id_63 ; give_act_reap; latency_task; check_ans;
	give_id_64 ; give_act_reap; latency_task; check_ans;
	give_id_65 ; give_act_reap; latency_task; check_ans;
	give_id_66 ; give_act_reap; latency_task; check_ans;
	give_id_67 ; give_act_reap; latency_task; check_ans;
	give_id_68 ; give_act_reap; latency_task; check_ans;
	give_id_69 ; give_act_reap; latency_task; check_ans;
	give_id_70 ; give_act_reap; latency_task; check_ans;
	give_id_71 ; give_act_reap; latency_task; check_ans;
	give_id_72 ; give_act_reap; latency_task; check_ans;
	give_id_73 ; give_act_reap; latency_task; check_ans;
	give_id_74 ; give_act_reap; latency_task; check_ans;
	give_id_75 ; give_act_reap; latency_task; check_ans;
	give_id_76 ; give_act_reap; latency_task; check_ans;
	give_id_77 ; give_act_reap; latency_task; check_ans;
	give_id_78 ; give_act_reap; latency_task; check_ans;
	give_id_79 ; give_act_reap; latency_task; check_ans;
	give_id_80 ; give_act_reap; latency_task; check_ans;
	give_id_81 ; give_act_reap; latency_task; check_ans;
	give_id_82 ; give_act_reap; latency_task; check_ans;
	give_id_83 ; give_act_reap; latency_task; check_ans;
	give_id_84 ; give_act_reap; latency_task; check_ans;
	give_id_85 ; give_act_reap; latency_task; check_ans;
	give_id_86 ; give_act_reap; latency_task; check_ans;
	give_id_87 ; give_act_reap; latency_task; check_ans;
	give_id_88 ; give_act_reap; latency_task; check_ans;
	give_id_89 ; give_act_reap; latency_task; check_ans;
	give_id_90 ; give_act_reap; latency_task; check_ans;
	give_id_91 ; give_act_reap; latency_task; check_ans;
	give_id_92 ; give_act_reap; latency_task; check_ans;
	give_id_93 ; give_act_reap; latency_task; check_ans;
	give_id_94 ; give_act_reap; latency_task; check_ans;
	give_id_95 ; give_act_reap; latency_task; check_ans;
	give_id_96 ; give_act_reap; latency_task; check_ans;
	give_id_97 ; give_act_reap; latency_task; check_ans;
	give_id_98 ; give_act_reap; latency_task; check_ans;
	give_id_99 ; give_act_reap; latency_task; check_ans;
	give_id_100; give_act_reap; latency_task; check_ans;
	give_id_101; give_act_reap; latency_task; check_ans;
	give_id_102; give_act_reap; latency_task; check_ans;
	give_id_103; give_act_reap; latency_task; check_ans;
	give_id_104; give_act_reap; latency_task; check_ans;
	give_id_105; give_act_reap; latency_task; check_ans;
	give_id_106; give_act_reap; latency_task; check_ans;
	give_id_107; give_act_reap; latency_task; check_ans;
	give_id_108; give_act_reap; latency_task; check_ans;
	give_id_109; give_act_reap; latency_task; check_ans;
	give_id_110; give_act_reap; latency_task; check_ans;
	give_id_111; give_act_reap; latency_task; check_ans;
	give_id_112; give_act_reap; latency_task; check_ans;
	give_id_113; give_act_reap; latency_task; check_ans;
	give_id_114; give_act_reap; latency_task; check_ans;
	give_id_115; give_act_reap; latency_task; check_ans;
	give_id_116; give_act_reap; latency_task; check_ans;
	give_id_117; give_act_reap; latency_task; check_ans;
	give_id_118; give_act_reap; latency_task; check_ans;
	give_id_119; give_act_reap; latency_task; check_ans;
	give_id_120; give_act_reap; latency_task; check_ans;
	give_id_121; give_act_reap; latency_task; check_ans;
	give_id_122; give_act_reap; latency_task; check_ans;
	give_id_123; give_act_reap; latency_task; check_ans;
	give_id_124; give_act_reap; latency_task; check_ans;
	give_id_125; give_act_reap; latency_task; check_ans;
	give_id_126; give_act_reap; latency_task; check_ans;
	give_id_127; give_act_reap; latency_task; check_ans;
	give_id_128; give_act_reap; latency_task; check_ans;
	give_id_129; give_act_reap; latency_task; check_ans;
	give_id_130; give_act_reap; latency_task; check_ans;
	give_id_131; give_act_reap; latency_task; check_ans;
	give_id_132; give_act_reap; latency_task; check_ans;
	give_id_133; give_act_reap; latency_task; check_ans;
	give_id_134; give_act_reap; latency_task; check_ans;
	give_id_135; give_act_reap; latency_task; check_ans;
	give_id_136; give_act_reap; latency_task; check_ans;
	give_id_137; give_act_reap; latency_task; check_ans;
	give_id_138; give_act_reap; latency_task; check_ans;
	give_id_139; give_act_reap; latency_task; check_ans;
	give_id_140; give_act_reap; latency_task; check_ans;
	give_id_141; give_act_reap; latency_task; check_ans;
	give_id_142; give_act_reap; latency_task; check_ans;
	give_id_143; give_act_reap; latency_task; check_ans;
	give_id_144; give_act_reap; latency_task; check_ans;
	give_id_145; give_act_reap; latency_task; check_ans;
	give_id_146; give_act_reap; latency_task; check_ans;
	give_id_147; give_act_reap; latency_task; check_ans;
	give_id_148; give_act_reap; latency_task; check_ans;
	give_id_149; give_act_reap; latency_task; check_ans;
	give_id_150; give_act_reap; latency_task; check_ans;
	give_id_151; give_act_reap; latency_task; check_ans;
	give_id_152; give_act_reap; latency_task; check_ans;
	give_id_153; give_act_reap; latency_task; check_ans;
	give_id_154; give_act_reap; latency_task; check_ans;
	give_id_155; give_act_reap; latency_task; check_ans;
	give_id_156; give_act_reap; latency_task; check_ans;
	give_id_157; give_act_reap; latency_task; check_ans;
	give_id_158; give_act_reap; latency_task; check_ans;
	give_id_159; give_act_reap; latency_task; check_ans;
	give_id_160; give_act_reap; latency_task; check_ans;
	give_id_161; give_act_reap; latency_task; check_ans;
	give_id_162; give_act_reap; latency_task; check_ans;
	give_id_163; give_act_reap; latency_task; check_ans;
	give_id_164; give_act_reap; latency_task; check_ans;
	give_id_165; give_act_reap; latency_task; check_ans;
	give_id_166; give_act_reap; latency_task; check_ans;
	give_id_167; give_act_reap; latency_task; check_ans;
	give_id_168; give_act_reap; latency_task; check_ans;
	give_id_169; give_act_reap; latency_task; check_ans;
	give_id_170; give_act_reap; latency_task; check_ans;
	give_id_171; give_act_reap; latency_task; check_ans;
	give_id_172; give_act_reap; latency_task; check_ans;
	give_id_173; give_act_reap; latency_task; check_ans;
	give_id_174; give_act_reap; latency_task; check_ans;
	give_id_175; give_act_reap; latency_task; check_ans;
	give_id_176; give_act_reap; latency_task; check_ans;
	give_id_177; give_act_reap; latency_task; check_ans;
	give_id_178; give_act_reap; latency_task; check_ans;
	give_id_179; give_act_reap; latency_task; check_ans;
	give_id_180; give_act_reap; latency_task; check_ans;
	give_id_181; give_act_reap; latency_task; check_ans;
	give_id_182; give_act_reap; latency_task; check_ans;
	give_id_183; give_act_reap; latency_task; check_ans;
	give_id_184; give_act_reap; latency_task; check_ans;
	give_id_185; give_act_reap; latency_task; check_ans;
	give_id_186; give_act_reap; latency_task; check_ans;
	give_id_187; give_act_reap; latency_task; check_ans;
	give_id_188; give_act_reap; latency_task; check_ans;
	give_id_189; give_act_reap; latency_task; check_ans;
	give_id_190; give_act_reap; latency_task; check_ans;
	give_id_191; give_act_reap; latency_task; check_ans;
	give_id_192; give_act_reap; latency_task; check_ans;
	give_id_193; give_act_reap; latency_task; check_ans;
	give_id_194; give_act_reap; latency_task; check_ans;
	give_id_195; give_act_reap; latency_task; check_ans;
	give_id_196; give_act_reap; latency_task; check_ans;
	give_id_197; give_act_reap; latency_task; check_ans;
	give_id_198; give_act_reap; latency_task; check_ans;
	give_id_199; give_act_reap; latency_task; check_ans;
	give_id_200; give_act_reap; latency_task; check_ans;
	give_id_201; give_act_reap; latency_task; check_ans;
	give_id_202; give_act_reap; latency_task; check_ans;
	give_id_203; give_act_reap; latency_task; check_ans;
	give_id_204; give_act_reap; latency_task; check_ans;
	give_id_205; give_act_reap; latency_task; check_ans;
	give_id_206; give_act_reap; latency_task; check_ans;
	give_id_207; give_act_reap; latency_task; check_ans;
	give_id_208; give_act_reap; latency_task; check_ans;
	give_id_209; give_act_reap; latency_task; check_ans;
	give_id_210; give_act_reap; latency_task; check_ans;
	give_id_211; give_act_reap; latency_task; check_ans;
	give_id_212; give_act_reap; latency_task; check_ans;
	give_id_213; give_act_reap; latency_task; check_ans;
	give_id_214; give_act_reap; latency_task; check_ans;
	give_id_215; give_act_reap; latency_task; check_ans;
	give_id_216; give_act_reap; latency_task; check_ans;
	give_id_217; give_act_reap; latency_task; check_ans;
	give_id_218; give_act_reap; latency_task; check_ans;
	give_id_219; give_act_reap; latency_task; check_ans;
	give_id_220; give_act_reap; latency_task; check_ans;
	give_id_221; give_act_reap; latency_task; check_ans;
	give_id_222; give_act_reap; latency_task; check_ans;
	give_id_223; give_act_reap; latency_task; check_ans;
	give_id_224; give_act_reap; latency_task; check_ans;
	give_id_225; give_act_reap; latency_task; check_ans;
	give_id_226; give_act_reap; latency_task; check_ans;
	give_id_227; give_act_reap; latency_task; check_ans;
	give_id_228; give_act_reap; latency_task; check_ans;
	give_id_229; give_act_reap; latency_task; check_ans;
	give_id_230; give_act_reap; latency_task; check_ans;
	give_id_231; give_act_reap; latency_task; check_ans;
	give_id_232; give_act_reap; latency_task; check_ans;
	give_id_233; give_act_reap; latency_task; check_ans;
	give_id_234; give_act_reap; latency_task; check_ans;
	give_id_235; give_act_reap; latency_task; check_ans;
	give_id_236; give_act_reap; latency_task; check_ans;
	give_id_237; give_act_reap; latency_task; check_ans;
	give_id_238; give_act_reap; latency_task; check_ans;
	give_id_239; give_act_reap; latency_task; check_ans;
	give_id_240; give_act_reap; latency_task; check_ans;
	give_id_241; give_act_reap; latency_task; check_ans;
	give_id_242; give_act_reap; latency_task; check_ans;
	give_id_243; give_act_reap; latency_task; check_ans;
	give_id_244; give_act_reap; latency_task; check_ans;
	give_id_245; give_act_reap; latency_task; check_ans;
	give_id_246; give_act_reap; latency_task; check_ans;
	give_id_247; give_act_reap; latency_task; check_ans;
	give_id_248; give_act_reap; latency_task; check_ans;
	give_id_249; give_act_reap; latency_task; check_ans;
	give_id_250; give_act_reap; latency_task; check_ans;
	give_id_251; give_act_reap; latency_task; check_ans;
	give_id_252; give_act_reap; latency_task; check_ans;
	give_id_253; give_act_reap; latency_task; check_ans;
	give_id_254; give_act_reap; latency_task; check_ans;
	// ID 4
	give_id_0  ; give_act_reap; latency_task; check_ans;
	give_id_1  ; give_act_reap; latency_task; check_ans;
	give_id_2  ; give_act_reap; latency_task; check_ans;
	give_id_3  ; give_act_reap; latency_task; check_ans;
	give_id_4  ; give_act_reap; latency_task; check_ans;
	give_id_5  ; give_act_reap; latency_task; check_ans;
	give_id_6  ; give_act_reap; latency_task; check_ans;
	give_id_7  ; give_act_reap; latency_task; check_ans;
	give_id_8  ; give_act_reap; latency_task; check_ans;
	give_id_9  ; give_act_reap; latency_task; check_ans;
	give_id_10 ; give_act_reap; latency_task; check_ans;
	give_id_11 ; give_act_reap; latency_task; check_ans;
	give_id_12 ; give_act_reap; latency_task; check_ans;
	give_id_13 ; give_act_reap; latency_task; check_ans;
	give_id_14 ; give_act_reap; latency_task; check_ans;
	give_id_15 ; give_act_reap; latency_task; check_ans;
	give_id_16 ; give_act_reap; latency_task; check_ans;
	give_id_17 ; give_act_reap; latency_task; check_ans;
	give_id_18 ; give_act_reap; latency_task; check_ans;
	give_id_19 ; give_act_reap; latency_task; check_ans;
	give_id_20 ; give_act_reap; latency_task; check_ans;
	give_id_21 ; give_act_reap; latency_task; check_ans;
	give_id_22 ; give_act_reap; latency_task; check_ans;
	give_id_23 ; give_act_reap; latency_task; check_ans;
	give_id_24 ; give_act_reap; latency_task; check_ans;
	give_id_25 ; give_act_reap; latency_task; check_ans;
	give_id_26 ; give_act_reap; latency_task; check_ans;
	give_id_27 ; give_act_reap; latency_task; check_ans;
	give_id_28 ; give_act_reap; latency_task; check_ans;
	give_id_29 ; give_act_reap; latency_task; check_ans;
	give_id_30 ; give_act_reap; latency_task; check_ans;
	give_id_31 ; give_act_reap; latency_task; check_ans;
	give_id_32 ; give_act_reap; latency_task; check_ans;
	give_id_33 ; give_act_reap; latency_task; check_ans;
	give_id_34 ; give_act_reap; latency_task; check_ans;
	give_id_35 ; give_act_reap; latency_task; check_ans;
	give_id_36 ; give_act_reap; latency_task; check_ans;
	give_id_37 ; give_act_reap; latency_task; check_ans;
	give_id_38 ; give_act_reap; latency_task; check_ans;
	give_id_39 ; give_act_reap; latency_task; check_ans;
	give_id_40 ; give_act_reap; latency_task; check_ans;
	give_id_41 ; give_act_reap; latency_task; check_ans;
	give_id_42 ; give_act_reap; latency_task; check_ans;
	give_id_43 ; give_act_reap; latency_task; check_ans;
	give_id_44 ; give_act_reap; latency_task; check_ans;
	give_id_45 ; give_act_reap; latency_task; check_ans;
	give_id_46 ; give_act_reap; latency_task; check_ans;
	give_id_47 ; give_act_reap; latency_task; check_ans;
	give_id_48 ; give_act_reap; latency_task; check_ans;
	give_id_49 ; give_act_reap; latency_task; check_ans;
	give_id_50 ; give_act_reap; latency_task; check_ans;
	give_id_51 ; give_act_reap; latency_task; check_ans;
	give_id_52 ; give_act_reap; latency_task; check_ans;
	give_id_53 ; give_act_reap; latency_task; check_ans;
	give_id_54 ; give_act_reap; latency_task; check_ans;
	give_id_55 ; give_act_reap; latency_task; check_ans;
	give_id_56 ; give_act_reap; latency_task; check_ans;
	give_id_57 ; give_act_reap; latency_task; check_ans;
	give_id_58 ; give_act_reap; latency_task; check_ans;
	give_id_59 ; give_act_reap; latency_task; check_ans;
	give_id_60 ; give_act_reap; latency_task; check_ans;
	give_id_61 ; give_act_reap; latency_task; check_ans;
	give_id_62 ; give_act_reap; latency_task; check_ans;
	give_id_63 ; give_act_reap; latency_task; check_ans;
	give_id_64 ; give_act_reap; latency_task; check_ans;
	give_id_65 ; give_act_reap; latency_task; check_ans;
	give_id_66 ; give_act_reap; latency_task; check_ans;
	give_id_67 ; give_act_reap; latency_task; check_ans;
	give_id_68 ; give_act_reap; latency_task; check_ans;
	give_id_69 ; give_act_reap; latency_task; check_ans;
	give_id_70 ; give_act_reap; latency_task; check_ans;
	give_id_71 ; give_act_reap; latency_task; check_ans;
	give_id_72 ; give_act_reap; latency_task; check_ans;
	give_id_73 ; give_act_reap; latency_task; check_ans;
	give_id_74 ; give_act_reap; latency_task; check_ans;
	give_id_75 ; give_act_reap; latency_task; check_ans;
	give_id_76 ; give_act_reap; latency_task; check_ans;
	give_id_77 ; give_act_reap; latency_task; check_ans;
	give_id_78 ; give_act_reap; latency_task; check_ans;
	give_id_79 ; give_act_reap; latency_task; check_ans;
	give_id_80 ; give_act_reap; latency_task; check_ans;
	give_id_81 ; give_act_reap; latency_task; check_ans;
	give_id_82 ; give_act_reap; latency_task; check_ans;
	give_id_83 ; give_act_reap; latency_task; check_ans;
	give_id_84 ; give_act_reap; latency_task; check_ans;
	give_id_85 ; give_act_reap; latency_task; check_ans;
	give_id_86 ; give_act_reap; latency_task; check_ans;
	give_id_87 ; give_act_reap; latency_task; check_ans;
	give_id_88 ; give_act_reap; latency_task; check_ans;
	give_id_89 ; give_act_reap; latency_task; check_ans;
	give_id_90 ; give_act_reap; latency_task; check_ans;
	give_id_91 ; give_act_reap; latency_task; check_ans;
	give_id_92 ; give_act_reap; latency_task; check_ans;
	give_id_93 ; give_act_reap; latency_task; check_ans;
	give_id_94 ; give_act_reap; latency_task; check_ans;
	give_id_95 ; give_act_reap; latency_task; check_ans;
	give_id_96 ; give_act_reap; latency_task; check_ans;
	give_id_97 ; give_act_reap; latency_task; check_ans;
	give_id_98 ; give_act_reap; latency_task; check_ans;
	give_id_99 ; give_act_reap; latency_task; check_ans;
	give_id_100; give_act_reap; latency_task; check_ans;
	give_id_101; give_act_reap; latency_task; check_ans;
	give_id_102; give_act_reap; latency_task; check_ans;
	give_id_103; give_act_reap; latency_task; check_ans;
	give_id_104; give_act_reap; latency_task; check_ans;
	give_id_105; give_act_reap; latency_task; check_ans;
	give_id_106; give_act_reap; latency_task; check_ans;
	give_id_107; give_act_reap; latency_task; check_ans;
	give_id_108; give_act_reap; latency_task; check_ans;
	give_id_109; give_act_reap; latency_task; check_ans;
	give_id_110; give_act_reap; latency_task; check_ans;
	give_id_111; give_act_reap; latency_task; check_ans;
	give_id_112; give_act_reap; latency_task; check_ans;
	give_id_113; give_act_reap; latency_task; check_ans;
	give_id_114; give_act_reap; latency_task; check_ans;
	give_id_115; give_act_reap; latency_task; check_ans;
	give_id_116; give_act_reap; latency_task; check_ans;
	give_id_117; give_act_reap; latency_task; check_ans;
	give_id_118; give_act_reap; latency_task; check_ans;
	give_id_119; give_act_reap; latency_task; check_ans;
	give_id_120; give_act_reap; latency_task; check_ans;
	give_id_121; give_act_reap; latency_task; check_ans;
	give_id_122; give_act_reap; latency_task; check_ans;
	give_id_123; give_act_reap; latency_task; check_ans;
	give_id_124; give_act_reap; latency_task; check_ans;
	give_id_125; give_act_reap; latency_task; check_ans;
	give_id_126; give_act_reap; latency_task; check_ans;
	give_id_127; give_act_reap; latency_task; check_ans;
	give_id_128; give_act_reap; latency_task; check_ans;
	give_id_129; give_act_reap; latency_task; check_ans;
	give_id_130; give_act_reap; latency_task; check_ans;
	give_id_131; give_act_reap; latency_task; check_ans;
	give_id_132; give_act_reap; latency_task; check_ans;
	give_id_133; give_act_reap; latency_task; check_ans;
	give_id_134; give_act_reap; latency_task; check_ans;
	give_id_135; give_act_reap; latency_task; check_ans;
	give_id_136; give_act_reap; latency_task; check_ans;
	give_id_137; give_act_reap; latency_task; check_ans;
	give_id_138; give_act_reap; latency_task; check_ans;
	give_id_139; give_act_reap; latency_task; check_ans;
	give_id_140; give_act_reap; latency_task; check_ans;
	give_id_141; give_act_reap; latency_task; check_ans;
	give_id_142; give_act_reap; latency_task; check_ans;
	give_id_143; give_act_reap; latency_task; check_ans;
	give_id_144; give_act_reap; latency_task; check_ans;
	give_id_145; give_act_reap; latency_task; check_ans;
	give_id_146; give_act_reap; latency_task; check_ans;
	give_id_147; give_act_reap; latency_task; check_ans;
	give_id_148; give_act_reap; latency_task; check_ans;
	give_id_149; give_act_reap; latency_task; check_ans;
	give_id_150; give_act_reap; latency_task; check_ans;
	give_id_151; give_act_reap; latency_task; check_ans;
	give_id_152; give_act_reap; latency_task; check_ans;
	give_id_153; give_act_reap; latency_task; check_ans;
	give_id_154; give_act_reap; latency_task; check_ans;
	give_id_155; give_act_reap; latency_task; check_ans;
	give_id_156; give_act_reap; latency_task; check_ans;
	give_id_157; give_act_reap; latency_task; check_ans;
	give_id_158; give_act_reap; latency_task; check_ans;
	give_id_159; give_act_reap; latency_task; check_ans;
	give_id_160; give_act_reap; latency_task; check_ans;
	give_id_161; give_act_reap; latency_task; check_ans;
	give_id_162; give_act_reap; latency_task; check_ans;
	give_id_163; give_act_reap; latency_task; check_ans;
	give_id_164; give_act_reap; latency_task; check_ans;
	give_id_165; give_act_reap; latency_task; check_ans;
	give_id_166; give_act_reap; latency_task; check_ans;
	give_id_167; give_act_reap; latency_task; check_ans;
	give_id_168; give_act_reap; latency_task; check_ans;
	give_id_169; give_act_reap; latency_task; check_ans;
	give_id_170; give_act_reap; latency_task; check_ans;
	give_id_171; give_act_reap; latency_task; check_ans;
	give_id_172; give_act_reap; latency_task; check_ans;
	give_id_173; give_act_reap; latency_task; check_ans;
	give_id_174; give_act_reap; latency_task; check_ans;
	give_id_175; give_act_reap; latency_task; check_ans;
	give_id_176; give_act_reap; latency_task; check_ans;
	give_id_177; give_act_reap; latency_task; check_ans;
	give_id_178; give_act_reap; latency_task; check_ans;
	give_id_179; give_act_reap; latency_task; check_ans;
	give_id_180; give_act_reap; latency_task; check_ans;
	give_id_181; give_act_reap; latency_task; check_ans;
	give_id_182; give_act_reap; latency_task; check_ans;
	give_id_183; give_act_reap; latency_task; check_ans;
	give_id_184; give_act_reap; latency_task; check_ans;
	give_id_185; give_act_reap; latency_task; check_ans;
	give_id_186; give_act_reap; latency_task; check_ans;
	give_id_187; give_act_reap; latency_task; check_ans;
	give_id_188; give_act_reap; latency_task; check_ans;
	give_id_189; give_act_reap; latency_task; check_ans;
	give_id_190; give_act_reap; latency_task; check_ans;
	give_id_191; give_act_reap; latency_task; check_ans;
	give_id_192; give_act_reap; latency_task; check_ans;
	give_id_193; give_act_reap; latency_task; check_ans;
	give_id_194; give_act_reap; latency_task; check_ans;
	give_id_195; give_act_reap; latency_task; check_ans;
	give_id_196; give_act_reap; latency_task; check_ans;
	give_id_197; give_act_reap; latency_task; check_ans;
	give_id_198; give_act_reap; latency_task; check_ans;
	give_id_199; give_act_reap; latency_task; check_ans;
	give_id_200; give_act_reap; latency_task; check_ans;
	give_id_201; give_act_reap; latency_task; check_ans;
	give_id_202; give_act_reap; latency_task; check_ans;
	give_id_203; give_act_reap; latency_task; check_ans;
	give_id_204; give_act_reap; latency_task; check_ans;
	give_id_205; give_act_reap; latency_task; check_ans;
	give_id_206; give_act_reap; latency_task; check_ans;
	give_id_207; give_act_reap; latency_task; check_ans;
	give_id_208; give_act_reap; latency_task; check_ans;
	give_id_209; give_act_reap; latency_task; check_ans;
	give_id_210; give_act_reap; latency_task; check_ans;
	give_id_211; give_act_reap; latency_task; check_ans;
	give_id_212; give_act_reap; latency_task; check_ans;
	give_id_213; give_act_reap; latency_task; check_ans;
	give_id_214; give_act_reap; latency_task; check_ans;
	give_id_215; give_act_reap; latency_task; check_ans;
	give_id_216; give_act_reap; latency_task; check_ans;
	give_id_217; give_act_reap; latency_task; check_ans;
	give_id_218; give_act_reap; latency_task; check_ans;
	give_id_219; give_act_reap; latency_task; check_ans;
	give_id_220; give_act_reap; latency_task; check_ans;
	give_id_221; give_act_reap; latency_task; check_ans;
	give_id_222; give_act_reap; latency_task; check_ans;
	give_id_223; give_act_reap; latency_task; check_ans;
	give_id_224; give_act_reap; latency_task; check_ans;
	give_id_225; give_act_reap; latency_task; check_ans;
	give_id_226; give_act_reap; latency_task; check_ans;
	give_id_227; give_act_reap; latency_task; check_ans;
	give_id_228; give_act_reap; latency_task; check_ans;
	give_id_229; give_act_reap; latency_task; check_ans;
	give_id_230; give_act_reap; latency_task; check_ans;
	give_id_231; give_act_reap; latency_task; check_ans;
	give_id_232; give_act_reap; latency_task; check_ans;
	give_id_233; give_act_reap; latency_task; check_ans;
	give_id_234; give_act_reap; latency_task; check_ans;
	give_id_235; give_act_reap; latency_task; check_ans;
	give_id_236; give_act_reap; latency_task; check_ans;
	give_id_237; give_act_reap; latency_task; check_ans;
	give_id_238; give_act_reap; latency_task; check_ans;
	give_id_239; give_act_reap; latency_task; check_ans;
	give_id_240; give_act_reap; latency_task; check_ans;
	give_id_241; give_act_reap; latency_task; check_ans;
	give_id_242; give_act_reap; latency_task; check_ans;
	give_id_243; give_act_reap; latency_task; check_ans;
	give_id_244; give_act_reap; latency_task; check_ans;
	give_id_245; give_act_reap; latency_task; check_ans;
	give_id_246; give_act_reap; latency_task; check_ans;
	give_id_247; give_act_reap; latency_task; check_ans;
	give_id_248; give_act_reap; latency_task; check_ans;
	give_id_249; give_act_reap; latency_task; check_ans;
	give_id_250; give_act_reap; latency_task; check_ans;
	give_id_251; give_act_reap; latency_task; check_ans;
	give_id_252; give_act_reap; latency_task; check_ans;
	give_id_253; give_act_reap; latency_task; check_ans;
	give_id_254; give_act_reap; latency_task; check_ans;
	// ID 5
	give_id_0  ; give_act_reap; latency_task; check_ans;
	give_id_1  ; give_act_reap; latency_task; check_ans;
	give_id_2  ; give_act_reap; latency_task; check_ans;
	give_id_3  ; give_act_reap; latency_task; check_ans;
	give_id_4  ; give_act_reap; latency_task; check_ans;
	give_id_5  ; give_act_reap; latency_task; check_ans;
	give_id_6  ; give_act_reap; latency_task; check_ans;
	give_id_7  ; give_act_reap; latency_task; check_ans;
	give_id_8  ; give_act_reap; latency_task; check_ans;
	give_id_9  ; give_act_reap; latency_task; check_ans;
	give_id_10 ; give_act_reap; latency_task; check_ans;
	give_id_11 ; give_act_reap; latency_task; check_ans;
	give_id_12 ; give_act_reap; latency_task; check_ans;
	give_id_13 ; give_act_reap; latency_task; check_ans;
	give_id_14 ; give_act_reap; latency_task; check_ans;
	give_id_15 ; give_act_reap; latency_task; check_ans;
	give_id_16 ; give_act_reap; latency_task; check_ans;
	give_id_17 ; give_act_reap; latency_task; check_ans;
	give_id_18 ; give_act_reap; latency_task; check_ans;
	give_id_19 ; give_act_reap; latency_task; check_ans;
	give_id_20 ; give_act_reap; latency_task; check_ans;
	give_id_21 ; give_act_reap; latency_task; check_ans;
	give_id_22 ; give_act_reap; latency_task; check_ans;
	give_id_23 ; give_act_reap; latency_task; check_ans;
	give_id_24 ; give_act_reap; latency_task; check_ans;
	give_id_25 ; give_act_reap; latency_task; check_ans;
	give_id_26 ; give_act_reap; latency_task; check_ans;
	give_id_27 ; give_act_reap; latency_task; check_ans;
	give_id_28 ; give_act_reap; latency_task; check_ans;
	give_id_29 ; give_act_reap; latency_task; check_ans;
	give_id_30 ; give_act_reap; latency_task; check_ans;
	give_id_31 ; give_act_reap; latency_task; check_ans;
	give_id_32 ; give_act_reap; latency_task; check_ans;
	give_id_33 ; give_act_reap; latency_task; check_ans;
	give_id_34 ; give_act_reap; latency_task; check_ans;
	give_id_35 ; give_act_reap; latency_task; check_ans;
	give_id_36 ; give_act_reap; latency_task; check_ans;
	give_id_37 ; give_act_reap; latency_task; check_ans;
	give_id_38 ; give_act_reap; latency_task; check_ans;
	give_id_39 ; give_act_reap; latency_task; check_ans;
	give_id_40 ; give_act_reap; latency_task; check_ans;
	give_id_41 ; give_act_reap; latency_task; check_ans;
	give_id_42 ; give_act_reap; latency_task; check_ans;
	give_id_43 ; give_act_reap; latency_task; check_ans;
	give_id_44 ; give_act_reap; latency_task; check_ans;
	give_id_45 ; give_act_reap; latency_task; check_ans;
	give_id_46 ; give_act_reap; latency_task; check_ans;
	give_id_47 ; give_act_reap; latency_task; check_ans;
	give_id_48 ; give_act_reap; latency_task; check_ans;
	give_id_49 ; give_act_reap; latency_task; check_ans;
	give_id_50 ; give_act_reap; latency_task; check_ans;
	give_id_51 ; give_act_reap; latency_task; check_ans;
	give_id_52 ; give_act_reap; latency_task; check_ans;
	give_id_53 ; give_act_reap; latency_task; check_ans;
	give_id_54 ; give_act_reap; latency_task; check_ans;
	give_id_55 ; give_act_reap; latency_task; check_ans;
	give_id_56 ; give_act_reap; latency_task; check_ans;
	give_id_57 ; give_act_reap; latency_task; check_ans;
	give_id_58 ; give_act_reap; latency_task; check_ans;
	give_id_59 ; give_act_reap; latency_task; check_ans;
	give_id_60 ; give_act_reap; latency_task; check_ans;
	give_id_61 ; give_act_reap; latency_task; check_ans;
	give_id_62 ; give_act_reap; latency_task; check_ans;
	give_id_63 ; give_act_reap; latency_task; check_ans;
	give_id_64 ; give_act_reap; latency_task; check_ans;
	give_id_65 ; give_act_reap; latency_task; check_ans;
	give_id_66 ; give_act_reap; latency_task; check_ans;
	give_id_67 ; give_act_reap; latency_task; check_ans;
	give_id_68 ; give_act_reap; latency_task; check_ans;
	give_id_69 ; give_act_reap; latency_task; check_ans;
	give_id_70 ; give_act_reap; latency_task; check_ans;
	give_id_71 ; give_act_reap; latency_task; check_ans;
	give_id_72 ; give_act_reap; latency_task; check_ans;
	give_id_73 ; give_act_reap; latency_task; check_ans;
	give_id_74 ; give_act_reap; latency_task; check_ans;
	give_id_75 ; give_act_reap; latency_task; check_ans;
	give_id_76 ; give_act_reap; latency_task; check_ans;
	give_id_77 ; give_act_reap; latency_task; check_ans;
	give_id_78 ; give_act_reap; latency_task; check_ans;
	give_id_79 ; give_act_reap; latency_task; check_ans;
	give_id_80 ; give_act_reap; latency_task; check_ans;
	give_id_81 ; give_act_reap; latency_task; check_ans;
	give_id_82 ; give_act_reap; latency_task; check_ans;
	give_id_83 ; give_act_reap; latency_task; check_ans;
	give_id_84 ; give_act_reap; latency_task; check_ans;
	give_id_85 ; give_act_reap; latency_task; check_ans;
	give_id_86 ; give_act_reap; latency_task; check_ans;
	give_id_87 ; give_act_reap; latency_task; check_ans;
	give_id_88 ; give_act_reap; latency_task; check_ans;
	give_id_89 ; give_act_reap; latency_task; check_ans;
	give_id_90 ; give_act_reap; latency_task; check_ans;
	give_id_91 ; give_act_reap; latency_task; check_ans;
	give_id_92 ; give_act_reap; latency_task; check_ans;
	give_id_93 ; give_act_reap; latency_task; check_ans;
	give_id_94 ; give_act_reap; latency_task; check_ans;
	give_id_95 ; give_act_reap; latency_task; check_ans;
	give_id_96 ; give_act_reap; latency_task; check_ans;
	give_id_97 ; give_act_reap; latency_task; check_ans;
	give_id_98 ; give_act_reap; latency_task; check_ans;
	give_id_99 ; give_act_reap; latency_task; check_ans;
	give_id_100; give_act_reap; latency_task; check_ans;
	give_id_101; give_act_reap; latency_task; check_ans;
	give_id_102; give_act_reap; latency_task; check_ans;
	give_id_103; give_act_reap; latency_task; check_ans;
	give_id_104; give_act_reap; latency_task; check_ans;
	give_id_105; give_act_reap; latency_task; check_ans;
	give_id_106; give_act_reap; latency_task; check_ans;
	give_id_107; give_act_reap; latency_task; check_ans;
	give_id_108; give_act_reap; latency_task; check_ans;
	give_id_109; give_act_reap; latency_task; check_ans;
	give_id_110; give_act_reap; latency_task; check_ans;
	give_id_111; give_act_reap; latency_task; check_ans;
	give_id_112; give_act_reap; latency_task; check_ans;
	give_id_113; give_act_reap; latency_task; check_ans;
	give_id_114; give_act_reap; latency_task; check_ans;
	give_id_115; give_act_reap; latency_task; check_ans;
	give_id_116; give_act_reap; latency_task; check_ans;
	give_id_117; give_act_reap; latency_task; check_ans;
	give_id_118; give_act_reap; latency_task; check_ans;
	give_id_119; give_act_reap; latency_task; check_ans;
	give_id_120; give_act_reap; latency_task; check_ans;
	give_id_121; give_act_reap; latency_task; check_ans;
	give_id_122; give_act_reap; latency_task; check_ans;
	give_id_123; give_act_reap; latency_task; check_ans;
	give_id_124; give_act_reap; latency_task; check_ans;
	give_id_125; give_act_reap; latency_task; check_ans;
	give_id_126; give_act_reap; latency_task; check_ans;
	give_id_127; give_act_reap; latency_task; check_ans;
	give_id_128; give_act_reap; latency_task; check_ans;
	give_id_129; give_act_reap; latency_task; check_ans;
	give_id_130; give_act_reap; latency_task; check_ans;
	give_id_131; give_act_reap; latency_task; check_ans;
	give_id_132; give_act_reap; latency_task; check_ans;
	give_id_133; give_act_reap; latency_task; check_ans;
	give_id_134; give_act_reap; latency_task; check_ans;
	give_id_135; give_act_reap; latency_task; check_ans;
	give_id_136; give_act_reap; latency_task; check_ans;
	give_id_137; give_act_reap; latency_task; check_ans;
	give_id_138; give_act_reap; latency_task; check_ans;
	give_id_139; give_act_reap; latency_task; check_ans;
	give_id_140; give_act_reap; latency_task; check_ans;
	give_id_141; give_act_reap; latency_task; check_ans;
	give_id_142; give_act_reap; latency_task; check_ans;
	give_id_143; give_act_reap; latency_task; check_ans;
	give_id_144; give_act_reap; latency_task; check_ans;
	give_id_145; give_act_reap; latency_task; check_ans;
	give_id_146; give_act_reap; latency_task; check_ans;
	give_id_147; give_act_reap; latency_task; check_ans;
	give_id_148; give_act_reap; latency_task; check_ans;
	give_id_149; give_act_reap; latency_task; check_ans;
	give_id_150; give_act_reap; latency_task; check_ans;
	give_id_151; give_act_reap; latency_task; check_ans;
	give_id_152; give_act_reap; latency_task; check_ans;
	give_id_153; give_act_reap; latency_task; check_ans;
	give_id_154; give_act_reap; latency_task; check_ans;
	give_id_155; give_act_reap; latency_task; check_ans;
	give_id_156; give_act_reap; latency_task; check_ans;
	give_id_157; give_act_reap; latency_task; check_ans;
	give_id_158; give_act_reap; latency_task; check_ans;
	give_id_159; give_act_reap; latency_task; check_ans;
	give_id_160; give_act_reap; latency_task; check_ans;
	give_id_161; give_act_reap; latency_task; check_ans;
	give_id_162; give_act_reap; latency_task; check_ans;
	give_id_163; give_act_reap; latency_task; check_ans;
	give_id_164; give_act_reap; latency_task; check_ans;
	give_id_165; give_act_reap; latency_task; check_ans;
	give_id_166; give_act_reap; latency_task; check_ans;
	give_id_167; give_act_reap; latency_task; check_ans;
	give_id_168; give_act_reap; latency_task; check_ans;
	give_id_169; give_act_reap; latency_task; check_ans;
	give_id_170; give_act_reap; latency_task; check_ans;
	give_id_171; give_act_reap; latency_task; check_ans;
	give_id_172; give_act_reap; latency_task; check_ans;
	give_id_173; give_act_reap; latency_task; check_ans;
	give_id_174; give_act_reap; latency_task; check_ans;
	give_id_175; give_act_reap; latency_task; check_ans;
	give_id_176; give_act_reap; latency_task; check_ans;
	give_id_177; give_act_reap; latency_task; check_ans;
	give_id_178; give_act_reap; latency_task; check_ans;
	give_id_179; give_act_reap; latency_task; check_ans;
	give_id_180; give_act_reap; latency_task; check_ans;
	give_id_181; give_act_reap; latency_task; check_ans;
	give_id_182; give_act_reap; latency_task; check_ans;
	give_id_183; give_act_reap; latency_task; check_ans;
	give_id_184; give_act_reap; latency_task; check_ans;
	give_id_185; give_act_reap; latency_task; check_ans;
	give_id_186; give_act_reap; latency_task; check_ans;
	give_id_187; give_act_reap; latency_task; check_ans;
	give_id_188; give_act_reap; latency_task; check_ans;
	give_id_189; give_act_reap; latency_task; check_ans;
	give_id_190; give_act_reap; latency_task; check_ans;
	give_id_191; give_act_reap; latency_task; check_ans;
	give_id_192; give_act_reap; latency_task; check_ans;
	give_id_193; give_act_reap; latency_task; check_ans;
	give_id_194; give_act_reap; latency_task; check_ans;
	give_id_195; give_act_reap; latency_task; check_ans;
	give_id_196; give_act_reap; latency_task; check_ans;
	give_id_197; give_act_reap; latency_task; check_ans;
	give_id_198; give_act_reap; latency_task; check_ans;
	give_id_199; give_act_reap; latency_task; check_ans;
	give_id_200; give_act_reap; latency_task; check_ans;
	give_id_201; give_act_reap; latency_task; check_ans;
	give_id_202; give_act_reap; latency_task; check_ans;
	give_id_203; give_act_reap; latency_task; check_ans;
	give_id_204; give_act_reap; latency_task; check_ans;
	give_id_205; give_act_reap; latency_task; check_ans;
	give_id_206; give_act_reap; latency_task; check_ans;
	give_id_207; give_act_reap; latency_task; check_ans;
	give_id_208; give_act_reap; latency_task; check_ans;
	give_id_209; give_act_reap; latency_task; check_ans;
	give_id_210; give_act_reap; latency_task; check_ans;
	give_id_211; give_act_reap; latency_task; check_ans;
	give_id_212; give_act_reap; latency_task; check_ans;
	give_id_213; give_act_reap; latency_task; check_ans;
	give_id_214; give_act_reap; latency_task; check_ans;
	give_id_215; give_act_reap; latency_task; check_ans;
	give_id_216; give_act_reap; latency_task; check_ans;
	give_id_217; give_act_reap; latency_task; check_ans;
	give_id_218; give_act_reap; latency_task; check_ans;
	give_id_219; give_act_reap; latency_task; check_ans;
	give_id_220; give_act_reap; latency_task; check_ans;
	give_id_221; give_act_reap; latency_task; check_ans;
	give_id_222; give_act_reap; latency_task; check_ans;
	give_id_223; give_act_reap; latency_task; check_ans;
	give_id_224; give_act_reap; latency_task; check_ans;
	give_id_225; give_act_reap; latency_task; check_ans;
	give_id_226; give_act_reap; latency_task; check_ans;
	give_id_227; give_act_reap; latency_task; check_ans;
	give_id_228; give_act_reap; latency_task; check_ans;
	give_id_229; give_act_reap; latency_task; check_ans;
	give_id_230; give_act_reap; latency_task; check_ans;
	give_id_231; give_act_reap; latency_task; check_ans;
	give_id_232; give_act_reap; latency_task; check_ans;
	give_id_233; give_act_reap; latency_task; check_ans;
	give_id_234; give_act_reap; latency_task; check_ans;
	give_id_235; give_act_reap; latency_task; check_ans;
	give_id_236; give_act_reap; latency_task; check_ans;
	give_id_237; give_act_reap; latency_task; check_ans;
	give_id_238; give_act_reap; latency_task; check_ans;
	give_id_239; give_act_reap; latency_task; check_ans;
	give_id_240; give_act_reap; latency_task; check_ans;
	give_id_241; give_act_reap; latency_task; check_ans;
	give_id_242; give_act_reap; latency_task; check_ans;
	give_id_243; give_act_reap; latency_task; check_ans;
	give_id_244; give_act_reap; latency_task; check_ans;
	give_id_245; give_act_reap; latency_task; check_ans;
	give_id_246; give_act_reap; latency_task; check_ans;
	give_id_247; give_act_reap; latency_task; check_ans;
	give_id_248; give_act_reap; latency_task; check_ans;
	give_id_249; give_act_reap; latency_task; check_ans;
	give_id_250; give_act_reap; latency_task; check_ans;
	give_id_251; give_act_reap; latency_task; check_ans;
	give_id_252; give_act_reap; latency_task; check_ans;
	give_id_253; give_act_reap; latency_task; check_ans;
	give_id_254; give_act_reap; latency_task; check_ans;
	// ID 6
	give_id_0  ; give_act_reap; latency_task; check_ans;
	give_id_1  ; give_act_reap; latency_task; check_ans;
	give_id_2  ; give_act_reap; latency_task; check_ans;
	give_id_3  ; give_act_reap; latency_task; check_ans;
	give_id_4  ; give_act_reap; latency_task; check_ans;
	give_id_5  ; give_act_reap; latency_task; check_ans;
	give_id_6  ; give_act_reap; latency_task; check_ans;
	give_id_7  ; give_act_reap; latency_task; check_ans;
	give_id_8  ; give_act_reap; latency_task; check_ans;
	give_id_9  ; give_act_reap; latency_task; check_ans;
	give_id_10 ; give_act_reap; latency_task; check_ans;
	give_id_11 ; give_act_reap; latency_task; check_ans;
	give_id_12 ; give_act_reap; latency_task; check_ans;
	give_id_13 ; give_act_reap; latency_task; check_ans;
	give_id_14 ; give_act_reap; latency_task; check_ans;
	give_id_15 ; give_act_reap; latency_task; check_ans;
	give_id_16 ; give_act_reap; latency_task; check_ans;
	give_id_17 ; give_act_reap; latency_task; check_ans;
	give_id_18 ; give_act_reap; latency_task; check_ans;
	give_id_19 ; give_act_reap; latency_task; check_ans;
	give_id_20 ; give_act_reap; latency_task; check_ans;
	give_id_21 ; give_act_reap; latency_task; check_ans;
	give_id_22 ; give_act_reap; latency_task; check_ans;
	give_id_23 ; give_act_reap; latency_task; check_ans;
	give_id_24 ; give_act_reap; latency_task; check_ans;
	give_id_25 ; give_act_reap; latency_task; check_ans;
	give_id_26 ; give_act_reap; latency_task; check_ans;
	give_id_27 ; give_act_reap; latency_task; check_ans;
	give_id_28 ; give_act_reap; latency_task; check_ans;
	give_id_29 ; give_act_reap; latency_task; check_ans;
	give_id_30 ; give_act_reap; latency_task; check_ans;
	give_id_31 ; give_act_reap; latency_task; check_ans;
	give_id_32 ; give_act_reap; latency_task; check_ans;
	give_id_33 ; give_act_reap; latency_task; check_ans;
	give_id_34 ; give_act_reap; latency_task; check_ans;
	give_id_35 ; give_act_reap; latency_task; check_ans;
	give_id_36 ; give_act_reap; latency_task; check_ans;
	give_id_37 ; give_act_reap; latency_task; check_ans;
	give_id_38 ; give_act_reap; latency_task; check_ans;
	give_id_39 ; give_act_reap; latency_task; check_ans;
	give_id_40 ; give_act_reap; latency_task; check_ans;
	give_id_41 ; give_act_reap; latency_task; check_ans;
	give_id_42 ; give_act_reap; latency_task; check_ans;
	give_id_43 ; give_act_reap; latency_task; check_ans;
	give_id_44 ; give_act_reap; latency_task; check_ans;
	give_id_45 ; give_act_reap; latency_task; check_ans;
	give_id_46 ; give_act_reap; latency_task; check_ans;
	give_id_47 ; give_act_reap; latency_task; check_ans;
	give_id_48 ; give_act_reap; latency_task; check_ans;
	give_id_49 ; give_act_reap; latency_task; check_ans;
	give_id_50 ; give_act_reap; latency_task; check_ans;
	give_id_51 ; give_act_reap; latency_task; check_ans;
	give_id_52 ; give_act_reap; latency_task; check_ans;
	give_id_53 ; give_act_reap; latency_task; check_ans;
	give_id_54 ; give_act_reap; latency_task; check_ans;
	give_id_55 ; give_act_reap; latency_task; check_ans;
	give_id_56 ; give_act_reap; latency_task; check_ans;
	give_id_57 ; give_act_reap; latency_task; check_ans;
	give_id_58 ; give_act_reap; latency_task; check_ans;
	give_id_59 ; give_act_reap; latency_task; check_ans;
	give_id_60 ; give_act_reap; latency_task; check_ans;
	give_id_61 ; give_act_reap; latency_task; check_ans;
	give_id_62 ; give_act_reap; latency_task; check_ans;
	give_id_63 ; give_act_reap; latency_task; check_ans;
	give_id_64 ; give_act_reap; latency_task; check_ans;
	give_id_65 ; give_act_reap; latency_task; check_ans;
	give_id_66 ; give_act_reap; latency_task; check_ans;
	give_id_67 ; give_act_reap; latency_task; check_ans;
	give_id_68 ; give_act_reap; latency_task; check_ans;
	give_id_69 ; give_act_reap; latency_task; check_ans;
	give_id_70 ; give_act_reap; latency_task; check_ans;
	give_id_71 ; give_act_reap; latency_task; check_ans;
	give_id_72 ; give_act_reap; latency_task; check_ans;
	give_id_73 ; give_act_reap; latency_task; check_ans;
	give_id_74 ; give_act_reap; latency_task; check_ans;
	give_id_75 ; give_act_reap; latency_task; check_ans;
	give_id_76 ; give_act_reap; latency_task; check_ans;
	give_id_77 ; give_act_reap; latency_task; check_ans;
	give_id_78 ; give_act_reap; latency_task; check_ans;
	give_id_79 ; give_act_reap; latency_task; check_ans;
	give_id_80 ; give_act_reap; latency_task; check_ans;
	give_id_81 ; give_act_reap; latency_task; check_ans;
	give_id_82 ; give_act_reap; latency_task; check_ans;
	give_id_83 ; give_act_reap; latency_task; check_ans;
	give_id_84 ; give_act_reap; latency_task; check_ans;
	give_id_85 ; give_act_reap; latency_task; check_ans;
	give_id_86 ; give_act_reap; latency_task; check_ans;
	give_id_87 ; give_act_reap; latency_task; check_ans;
	give_id_88 ; give_act_reap; latency_task; check_ans;
	give_id_89 ; give_act_reap; latency_task; check_ans;
	give_id_90 ; give_act_reap; latency_task; check_ans;
	give_id_91 ; give_act_reap; latency_task; check_ans;
	give_id_92 ; give_act_reap; latency_task; check_ans;
	give_id_93 ; give_act_reap; latency_task; check_ans;
	give_id_94 ; give_act_reap; latency_task; check_ans;
	give_id_95 ; give_act_reap; latency_task; check_ans;
	give_id_96 ; give_act_reap; latency_task; check_ans;
	give_id_97 ; give_act_reap; latency_task; check_ans;
	give_id_98 ; give_act_reap; latency_task; check_ans;
	give_id_99 ; give_act_reap; latency_task; check_ans;
	give_id_100; give_act_reap; latency_task; check_ans;
	give_id_101; give_act_reap; latency_task; check_ans;
	give_id_102; give_act_reap; latency_task; check_ans;
	give_id_103; give_act_reap; latency_task; check_ans;
	give_id_104; give_act_reap; latency_task; check_ans;
	give_id_105; give_act_reap; latency_task; check_ans;
	give_id_106; give_act_reap; latency_task; check_ans;
	give_id_107; give_act_reap; latency_task; check_ans;
	give_id_108; give_act_reap; latency_task; check_ans;
	give_id_109; give_act_reap; latency_task; check_ans;
	give_id_110; give_act_reap; latency_task; check_ans;
	give_id_111; give_act_reap; latency_task; check_ans;
	give_id_112; give_act_reap; latency_task; check_ans;
	give_id_113; give_act_reap; latency_task; check_ans;
	give_id_114; give_act_reap; latency_task; check_ans;
	give_id_115; give_act_reap; latency_task; check_ans;
	give_id_116; give_act_reap; latency_task; check_ans;
	give_id_117; give_act_reap; latency_task; check_ans;
	give_id_118; give_act_reap; latency_task; check_ans;
	give_id_119; give_act_reap; latency_task; check_ans;
	give_id_120; give_act_reap; latency_task; check_ans;
	give_id_121; give_act_reap; latency_task; check_ans;
	give_id_122; give_act_reap; latency_task; check_ans;
	give_id_123; give_act_reap; latency_task; check_ans;
	give_id_124; give_act_reap; latency_task; check_ans;
	give_id_125; give_act_reap; latency_task; check_ans;
	give_id_126; give_act_reap; latency_task; check_ans;
	give_id_127; give_act_reap; latency_task; check_ans;
	give_id_128; give_act_reap; latency_task; check_ans;
	give_id_129; give_act_reap; latency_task; check_ans;
	give_id_130; give_act_reap; latency_task; check_ans;
	give_id_131; give_act_reap; latency_task; check_ans;
	give_id_132; give_act_reap; latency_task; check_ans;
	give_id_133; give_act_reap; latency_task; check_ans;
	give_id_134; give_act_reap; latency_task; check_ans;
	give_id_135; give_act_reap; latency_task; check_ans;
	give_id_136; give_act_reap; latency_task; check_ans;
	give_id_137; give_act_reap; latency_task; check_ans;
	give_id_138; give_act_reap; latency_task; check_ans;
	give_id_139; give_act_reap; latency_task; check_ans;
	give_id_140; give_act_reap; latency_task; check_ans;
	give_id_141; give_act_reap; latency_task; check_ans;
	give_id_142; give_act_reap; latency_task; check_ans;
	give_id_143; give_act_reap; latency_task; check_ans;
	give_id_144; give_act_reap; latency_task; check_ans;
	give_id_145; give_act_reap; latency_task; check_ans;
	give_id_146; give_act_reap; latency_task; check_ans;
	give_id_147; give_act_reap; latency_task; check_ans;
	give_id_148; give_act_reap; latency_task; check_ans;
	give_id_149; give_act_reap; latency_task; check_ans;
	give_id_150; give_act_reap; latency_task; check_ans;
	give_id_151; give_act_reap; latency_task; check_ans;
	give_id_152; give_act_reap; latency_task; check_ans;
	give_id_153; give_act_reap; latency_task; check_ans;
	give_id_154; give_act_reap; latency_task; check_ans;
	give_id_155; give_act_reap; latency_task; check_ans;
	give_id_156; give_act_reap; latency_task; check_ans;
	give_id_157; give_act_reap; latency_task; check_ans;
	give_id_158; give_act_reap; latency_task; check_ans;
	give_id_159; give_act_reap; latency_task; check_ans;
	give_id_160; give_act_reap; latency_task; check_ans;
	give_id_161; give_act_reap; latency_task; check_ans;
	give_id_162; give_act_reap; latency_task; check_ans;
	give_id_163; give_act_reap; latency_task; check_ans;
	give_id_164; give_act_reap; latency_task; check_ans;
	give_id_165; give_act_reap; latency_task; check_ans;
	give_id_166; give_act_reap; latency_task; check_ans;
	give_id_167; give_act_reap; latency_task; check_ans;
	give_id_168; give_act_reap; latency_task; check_ans;
	give_id_169; give_act_reap; latency_task; check_ans;
	give_id_170; give_act_reap; latency_task; check_ans;
	give_id_171; give_act_reap; latency_task; check_ans;
	give_id_172; give_act_reap; latency_task; check_ans;
	give_id_173; give_act_reap; latency_task; check_ans;
	give_id_174; give_act_reap; latency_task; check_ans;
	give_id_175; give_act_reap; latency_task; check_ans;
	give_id_176; give_act_reap; latency_task; check_ans;
	give_id_177; give_act_reap; latency_task; check_ans;
	give_id_178; give_act_reap; latency_task; check_ans;
	give_id_179; give_act_reap; latency_task; check_ans;
	give_id_180; give_act_reap; latency_task; check_ans;
	give_id_181; give_act_reap; latency_task; check_ans;
	give_id_182; give_act_reap; latency_task; check_ans;
	give_id_183; give_act_reap; latency_task; check_ans;
	give_id_184; give_act_reap; latency_task; check_ans;
	give_id_185; give_act_reap; latency_task; check_ans;
	give_id_186; give_act_reap; latency_task; check_ans;
	give_id_187; give_act_reap; latency_task; check_ans;
	give_id_188; give_act_reap; latency_task; check_ans;
	give_id_189; give_act_reap; latency_task; check_ans;
	give_id_190; give_act_reap; latency_task; check_ans;
	give_id_191; give_act_reap; latency_task; check_ans;
	give_id_192; give_act_reap; latency_task; check_ans;
	give_id_193; give_act_reap; latency_task; check_ans;
	give_id_194; give_act_reap; latency_task; check_ans;
	give_id_195; give_act_reap; latency_task; check_ans;
	give_id_196; give_act_reap; latency_task; check_ans;
	give_id_197; give_act_reap; latency_task; check_ans;
	give_id_198; give_act_reap; latency_task; check_ans;
	give_id_199; give_act_reap; latency_task; check_ans;
	give_id_200; give_act_reap; latency_task; check_ans;
	give_id_201; give_act_reap; latency_task; check_ans;
	give_id_202; give_act_reap; latency_task; check_ans;
	give_id_203; give_act_reap; latency_task; check_ans;
	give_id_204; give_act_reap; latency_task; check_ans;
	give_id_205; give_act_reap; latency_task; check_ans;
	give_id_206; give_act_reap; latency_task; check_ans;
	give_id_207; give_act_reap; latency_task; check_ans;
	give_id_208; give_act_reap; latency_task; check_ans;
	give_id_209; give_act_reap; latency_task; check_ans;
	give_id_210; give_act_reap; latency_task; check_ans;
	give_id_211; give_act_reap; latency_task; check_ans;
	give_id_212; give_act_reap; latency_task; check_ans;
	give_id_213; give_act_reap; latency_task; check_ans;
	give_id_214; give_act_reap; latency_task; check_ans;
	give_id_215; give_act_reap; latency_task; check_ans;
	give_id_216; give_act_reap; latency_task; check_ans;
	give_id_217; give_act_reap; latency_task; check_ans;
	give_id_218; give_act_reap; latency_task; check_ans;
	give_id_219; give_act_reap; latency_task; check_ans;
	give_id_220; give_act_reap; latency_task; check_ans;
	give_id_221; give_act_reap; latency_task; check_ans;
	give_id_222; give_act_reap; latency_task; check_ans;
	give_id_223; give_act_reap; latency_task; check_ans;
	give_id_224; give_act_reap; latency_task; check_ans;
	give_id_225; give_act_reap; latency_task; check_ans;
	give_id_226; give_act_reap; latency_task; check_ans;
	give_id_227; give_act_reap; latency_task; check_ans;
	give_id_228; give_act_reap; latency_task; check_ans;
	give_id_229; give_act_reap; latency_task; check_ans;
	give_id_230; give_act_reap; latency_task; check_ans;
	give_id_231; give_act_reap; latency_task; check_ans;
	give_id_232; give_act_reap; latency_task; check_ans;
	give_id_233; give_act_reap; latency_task; check_ans;
	give_id_234; give_act_reap; latency_task; check_ans;
	give_id_235; give_act_reap; latency_task; check_ans;
	give_id_236; give_act_reap; latency_task; check_ans;
	give_id_237; give_act_reap; latency_task; check_ans;
	give_id_238; give_act_reap; latency_task; check_ans;
	give_id_239; give_act_reap; latency_task; check_ans;
	give_id_240; give_act_reap; latency_task; check_ans;
	give_id_241; give_act_reap; latency_task; check_ans;
	give_id_242; give_act_reap; latency_task; check_ans;
	give_id_243; give_act_reap; latency_task; check_ans;
	give_id_244; give_act_reap; latency_task; check_ans;
	give_id_245; give_act_reap; latency_task; check_ans;
	give_id_246; give_act_reap; latency_task; check_ans;
	give_id_247; give_act_reap; latency_task; check_ans;
	give_id_248; give_act_reap; latency_task; check_ans;
	give_id_249; give_act_reap; latency_task; check_ans;
	give_id_250; give_act_reap; latency_task; check_ans;
	give_id_251; give_act_reap; latency_task; check_ans;
	give_id_252; give_act_reap; latency_task; check_ans;
	give_id_253; give_act_reap; latency_task; check_ans;
	give_id_254; give_act_reap; latency_task; check_ans;
	// ID 7
	give_id_0  ; give_act_reap; latency_task; check_ans;
	give_id_1  ; give_act_reap; latency_task; check_ans;
	give_id_2  ; give_act_reap; latency_task; check_ans;
	give_id_3  ; give_act_reap; latency_task; check_ans;
	give_id_4  ; give_act_reap; latency_task; check_ans;
	give_id_5  ; give_act_reap; latency_task; check_ans;
	give_id_6  ; give_act_reap; latency_task; check_ans;
	give_id_7  ; give_act_reap; latency_task; check_ans;
	give_id_8  ; give_act_reap; latency_task; check_ans;
	give_id_9  ; give_act_reap; latency_task; check_ans;
	give_id_10 ; give_act_reap; latency_task; check_ans;
	give_id_11 ; give_act_reap; latency_task; check_ans;
	give_id_12 ; give_act_reap; latency_task; check_ans;
	give_id_13 ; give_act_reap; latency_task; check_ans;
	give_id_14 ; give_act_reap; latency_task; check_ans;
	give_id_15 ; give_act_reap; latency_task; check_ans;
	give_id_16 ; give_act_reap; latency_task; check_ans;
	give_id_17 ; give_act_reap; latency_task; check_ans;
	give_id_18 ; give_act_reap; latency_task; check_ans;
	give_id_19 ; give_act_reap; latency_task; check_ans;
	give_id_20 ; give_act_reap; latency_task; check_ans;
	give_id_21 ; give_act_reap; latency_task; check_ans;
	give_id_22 ; give_act_reap; latency_task; check_ans;
	give_id_23 ; give_act_reap; latency_task; check_ans;
	give_id_24 ; give_act_reap; latency_task; check_ans;
	give_id_25 ; give_act_reap; latency_task; check_ans;
	give_id_26 ; give_act_reap; latency_task; check_ans;
	give_id_27 ; give_act_reap; latency_task; check_ans;
	give_id_28 ; give_act_reap; latency_task; check_ans;
	give_id_29 ; give_act_reap; latency_task; check_ans;
	give_id_30 ; give_act_reap; latency_task; check_ans;
	give_id_31 ; give_act_reap; latency_task; check_ans;
	give_id_32 ; give_act_reap; latency_task; check_ans;
	give_id_33 ; give_act_reap; latency_task; check_ans;
	give_id_34 ; give_act_reap; latency_task; check_ans;
	give_id_35 ; give_act_reap; latency_task; check_ans;
	give_id_36 ; give_act_reap; latency_task; check_ans;
	give_id_37 ; give_act_reap; latency_task; check_ans;
	give_id_38 ; give_act_reap; latency_task; check_ans;
	give_id_39 ; give_act_reap; latency_task; check_ans;
	give_id_40 ; give_act_reap; latency_task; check_ans;
	give_id_41 ; give_act_reap; latency_task; check_ans;
	give_id_42 ; give_act_reap; latency_task; check_ans;
	give_id_43 ; give_act_reap; latency_task; check_ans;
	give_id_44 ; give_act_reap; latency_task; check_ans;
	give_id_45 ; give_act_reap; latency_task; check_ans;
	give_id_46 ; give_act_reap; latency_task; check_ans;
	give_id_47 ; give_act_reap; latency_task; check_ans;
	give_id_48 ; give_act_reap; latency_task; check_ans;
	give_id_49 ; give_act_reap; latency_task; check_ans;
	give_id_50 ; give_act_reap; latency_task; check_ans;
	give_id_51 ; give_act_reap; latency_task; check_ans;
	give_id_52 ; give_act_reap; latency_task; check_ans;
	give_id_53 ; give_act_reap; latency_task; check_ans;
	give_id_54 ; give_act_reap; latency_task; check_ans;
	give_id_55 ; give_act_reap; latency_task; check_ans;
	give_id_56 ; give_act_reap; latency_task; check_ans;
	give_id_57 ; give_act_reap; latency_task; check_ans;
	give_id_58 ; give_act_reap; latency_task; check_ans;
	give_id_59 ; give_act_reap; latency_task; check_ans;
	give_id_60 ; give_act_reap; latency_task; check_ans;
	give_id_61 ; give_act_reap; latency_task; check_ans;
	give_id_62 ; give_act_reap; latency_task; check_ans;
	give_id_63 ; give_act_reap; latency_task; check_ans;
	give_id_64 ; give_act_reap; latency_task; check_ans;
	give_id_65 ; give_act_reap; latency_task; check_ans;
	give_id_66 ; give_act_reap; latency_task; check_ans;
	give_id_67 ; give_act_reap; latency_task; check_ans;
	give_id_68 ; give_act_reap; latency_task; check_ans;
	give_id_69 ; give_act_reap; latency_task; check_ans;
	give_id_70 ; give_act_reap; latency_task; check_ans;
	give_id_71 ; give_act_reap; latency_task; check_ans;
	give_id_72 ; give_act_reap; latency_task; check_ans;
	give_id_73 ; give_act_reap; latency_task; check_ans;
	give_id_74 ; give_act_reap; latency_task; check_ans;
	give_id_75 ; give_act_reap; latency_task; check_ans;
	give_id_76 ; give_act_reap; latency_task; check_ans;
	give_id_77 ; give_act_reap; latency_task; check_ans;
	give_id_78 ; give_act_reap; latency_task; check_ans;
	give_id_79 ; give_act_reap; latency_task; check_ans;
	give_id_80 ; give_act_reap; latency_task; check_ans;
	give_id_81 ; give_act_reap; latency_task; check_ans;
	give_id_82 ; give_act_reap; latency_task; check_ans;
	give_id_83 ; give_act_reap; latency_task; check_ans;
	give_id_84 ; give_act_reap; latency_task; check_ans;
	give_id_85 ; give_act_reap; latency_task; check_ans;
	give_id_86 ; give_act_reap; latency_task; check_ans;
	give_id_87 ; give_act_reap; latency_task; check_ans;
	give_id_88 ; give_act_reap; latency_task; check_ans;
	give_id_89 ; give_act_reap; latency_task; check_ans;
	give_id_90 ; give_act_reap; latency_task; check_ans;
	give_id_91 ; give_act_reap; latency_task; check_ans;
	give_id_92 ; give_act_reap; latency_task; check_ans;
	give_id_93 ; give_act_reap; latency_task; check_ans;
	give_id_94 ; give_act_reap; latency_task; check_ans;
	give_id_95 ; give_act_reap; latency_task; check_ans;
	give_id_96 ; give_act_reap; latency_task; check_ans;
	give_id_97 ; give_act_reap; latency_task; check_ans;
	give_id_98 ; give_act_reap; latency_task; check_ans;
	give_id_99 ; give_act_reap; latency_task; check_ans;
	give_id_100; give_act_reap; latency_task; check_ans;
	give_id_101; give_act_reap; latency_task; check_ans;
	give_id_102; give_act_reap; latency_task; check_ans;
	give_id_103; give_act_reap; latency_task; check_ans;
	give_id_104; give_act_reap; latency_task; check_ans;
	give_id_105; give_act_reap; latency_task; check_ans;
	give_id_106; give_act_reap; latency_task; check_ans;
	give_id_107; give_act_reap; latency_task; check_ans;
	give_id_108; give_act_reap; latency_task; check_ans;
	give_id_109; give_act_reap; latency_task; check_ans;
	give_id_110; give_act_reap; latency_task; check_ans;
	give_id_111; give_act_reap; latency_task; check_ans;
	give_id_112; give_act_reap; latency_task; check_ans;
	give_id_113; give_act_reap; latency_task; check_ans;
	give_id_114; give_act_reap; latency_task; check_ans;
	give_id_115; give_act_reap; latency_task; check_ans;
	give_id_116; give_act_reap; latency_task; check_ans;
	give_id_117; give_act_reap; latency_task; check_ans;
	give_id_118; give_act_reap; latency_task; check_ans;
	give_id_119; give_act_reap; latency_task; check_ans;
	give_id_120; give_act_reap; latency_task; check_ans;
	give_id_121; give_act_reap; latency_task; check_ans;
	give_id_122; give_act_reap; latency_task; check_ans;
	give_id_123; give_act_reap; latency_task; check_ans;
	give_id_124; give_act_reap; latency_task; check_ans;
	give_id_125; give_act_reap; latency_task; check_ans;
	give_id_126; give_act_reap; latency_task; check_ans;
	give_id_127; give_act_reap; latency_task; check_ans;
	give_id_128; give_act_reap; latency_task; check_ans;
	give_id_129; give_act_reap; latency_task; check_ans;
	give_id_130; give_act_reap; latency_task; check_ans;
	give_id_131; give_act_reap; latency_task; check_ans;
	give_id_132; give_act_reap; latency_task; check_ans;
	give_id_133; give_act_reap; latency_task; check_ans;
	give_id_134; give_act_reap; latency_task; check_ans;
	give_id_135; give_act_reap; latency_task; check_ans;
	give_id_136; give_act_reap; latency_task; check_ans;
	give_id_137; give_act_reap; latency_task; check_ans;
	give_id_138; give_act_reap; latency_task; check_ans;
	give_id_139; give_act_reap; latency_task; check_ans;
	give_id_140; give_act_reap; latency_task; check_ans;
	give_id_141; give_act_reap; latency_task; check_ans;
	give_id_142; give_act_reap; latency_task; check_ans;
	give_id_143; give_act_reap; latency_task; check_ans;
	give_id_144; give_act_reap; latency_task; check_ans;
	give_id_145; give_act_reap; latency_task; check_ans;
	give_id_146; give_act_reap; latency_task; check_ans;
	give_id_147; give_act_reap; latency_task; check_ans;
	give_id_148; give_act_reap; latency_task; check_ans;
	give_id_149; give_act_reap; latency_task; check_ans;
	give_id_150; give_act_reap; latency_task; check_ans;
	give_id_151; give_act_reap; latency_task; check_ans;
	give_id_152; give_act_reap; latency_task; check_ans;
	give_id_153; give_act_reap; latency_task; check_ans;
	give_id_154; give_act_reap; latency_task; check_ans;
	give_id_155; give_act_reap; latency_task; check_ans;
	give_id_156; give_act_reap; latency_task; check_ans;
	give_id_157; give_act_reap; latency_task; check_ans;
	give_id_158; give_act_reap; latency_task; check_ans;
	give_id_159; give_act_reap; latency_task; check_ans;
	give_id_160; give_act_reap; latency_task; check_ans;
	give_id_161; give_act_reap; latency_task; check_ans;
	give_id_162; give_act_reap; latency_task; check_ans;
	give_id_163; give_act_reap; latency_task; check_ans;
	give_id_164; give_act_reap; latency_task; check_ans;
	give_id_165; give_act_reap; latency_task; check_ans;
	give_id_166; give_act_reap; latency_task; check_ans;
	give_id_167; give_act_reap; latency_task; check_ans;
	give_id_168; give_act_reap; latency_task; check_ans;
	give_id_169; give_act_reap; latency_task; check_ans;
	give_id_170; give_act_reap; latency_task; check_ans;
	give_id_171; give_act_reap; latency_task; check_ans;
	give_id_172; give_act_reap; latency_task; check_ans;
	give_id_173; give_act_reap; latency_task; check_ans;
	give_id_174; give_act_reap; latency_task; check_ans;
	give_id_175; give_act_reap; latency_task; check_ans;
	give_id_176; give_act_reap; latency_task; check_ans;
	give_id_177; give_act_reap; latency_task; check_ans;
	give_id_178; give_act_reap; latency_task; check_ans;
	give_id_179; give_act_reap; latency_task; check_ans;
	give_id_180; give_act_reap; latency_task; check_ans;
	give_id_181; give_act_reap; latency_task; check_ans;
	give_id_182; give_act_reap; latency_task; check_ans;
	give_id_183; give_act_reap; latency_task; check_ans;
	give_id_184; give_act_reap; latency_task; check_ans;
	give_id_185; give_act_reap; latency_task; check_ans;
	give_id_186; give_act_reap; latency_task; check_ans;
	give_id_187; give_act_reap; latency_task; check_ans;
	give_id_188; give_act_reap; latency_task; check_ans;
	give_id_189; give_act_reap; latency_task; check_ans;
	give_id_190; give_act_reap; latency_task; check_ans;
	give_id_191; give_act_reap; latency_task; check_ans;
	give_id_192; give_act_reap; latency_task; check_ans;
	give_id_193; give_act_reap; latency_task; check_ans;
	give_id_194; give_act_reap; latency_task; check_ans;
	give_id_195; give_act_reap; latency_task; check_ans;
	give_id_196; give_act_reap; latency_task; check_ans;
	give_id_197; give_act_reap; latency_task; check_ans;
	give_id_198; give_act_reap; latency_task; check_ans;
	give_id_199; give_act_reap; latency_task; check_ans;
	give_id_200; give_act_reap; latency_task; check_ans;
	give_id_201; give_act_reap; latency_task; check_ans;
	give_id_202; give_act_reap; latency_task; check_ans;
	give_id_203; give_act_reap; latency_task; check_ans;
	give_id_204; give_act_reap; latency_task; check_ans;
	give_id_205; give_act_reap; latency_task; check_ans;
	give_id_206; give_act_reap; latency_task; check_ans;
	give_id_207; give_act_reap; latency_task; check_ans;
	give_id_208; give_act_reap; latency_task; check_ans;
	give_id_209; give_act_reap; latency_task; check_ans;
	give_id_210; give_act_reap; latency_task; check_ans;
	give_id_211; give_act_reap; latency_task; check_ans;
	give_id_212; give_act_reap; latency_task; check_ans;
	give_id_213; give_act_reap; latency_task; check_ans;
	give_id_214; give_act_reap; latency_task; check_ans;
	give_id_215; give_act_reap; latency_task; check_ans;
	give_id_216; give_act_reap; latency_task; check_ans;
	give_id_217; give_act_reap; latency_task; check_ans;
	give_id_218; give_act_reap; latency_task; check_ans;
	give_id_219; give_act_reap; latency_task; check_ans;
	give_id_220; give_act_reap; latency_task; check_ans;
	give_id_221; give_act_reap; latency_task; check_ans;
	give_id_222; give_act_reap; latency_task; check_ans;
	give_id_223; give_act_reap; latency_task; check_ans;
	give_id_224; give_act_reap; latency_task; check_ans;
	give_id_225; give_act_reap; latency_task; check_ans;
	give_id_226; give_act_reap; latency_task; check_ans;
	give_id_227; give_act_reap; latency_task; check_ans;
	give_id_228; give_act_reap; latency_task; check_ans;
	give_id_229; give_act_reap; latency_task; check_ans;
	give_id_230; give_act_reap; latency_task; check_ans;
	give_id_231; give_act_reap; latency_task; check_ans;
	give_id_232; give_act_reap; latency_task; check_ans;
	give_id_233; give_act_reap; latency_task; check_ans;
	give_id_234; give_act_reap; latency_task; check_ans;
	give_id_235; give_act_reap; latency_task; check_ans;
	give_id_236; give_act_reap; latency_task; check_ans;
	give_id_237; give_act_reap; latency_task; check_ans;
	give_id_238; give_act_reap; latency_task; check_ans;
	give_id_239; give_act_reap; latency_task; check_ans;
	give_id_240; give_act_reap; latency_task; check_ans;
	give_id_241; give_act_reap; latency_task; check_ans;
	give_id_242; give_act_reap; latency_task; check_ans;
	give_id_243; give_act_reap; latency_task; check_ans;
	give_id_244; give_act_reap; latency_task; check_ans;
	give_id_245; give_act_reap; latency_task; check_ans;
	give_id_246; give_act_reap; latency_task; check_ans;
	give_id_247; give_act_reap; latency_task; check_ans;
	give_id_248; give_act_reap; latency_task; check_ans;
	give_id_249; give_act_reap; latency_task; check_ans;
	give_id_250; give_act_reap; latency_task; check_ans;
	give_id_251; give_act_reap; latency_task; check_ans;
	give_id_252; give_act_reap; latency_task; check_ans;
	give_id_253; give_act_reap; latency_task; check_ans;
	give_id_254; give_act_reap; latency_task; check_ans;
	// ID 8
	give_id_0  ; give_act_reap; latency_task; check_ans;
	give_id_1  ; give_act_reap; latency_task; check_ans;
	give_id_2  ; give_act_reap; latency_task; check_ans;
	give_id_3  ; give_act_reap; latency_task; check_ans;
	give_id_4  ; give_act_reap; latency_task; check_ans;
	give_id_5  ; give_act_reap; latency_task; check_ans;
	give_id_6  ; give_act_reap; latency_task; check_ans;
	give_id_7  ; give_act_reap; latency_task; check_ans;
	give_id_8  ; give_act_reap; latency_task; check_ans;
	give_id_9  ; give_act_reap; latency_task; check_ans;
	give_id_10 ; give_act_reap; latency_task; check_ans;
	give_id_11 ; give_act_reap; latency_task; check_ans;
	give_id_12 ; give_act_reap; latency_task; check_ans;
	give_id_13 ; give_act_reap; latency_task; check_ans;
	give_id_14 ; give_act_reap; latency_task; check_ans;
	give_id_15 ; give_act_reap; latency_task; check_ans;
	give_id_16 ; give_act_reap; latency_task; check_ans;
	give_id_17 ; give_act_reap; latency_task; check_ans;
	give_id_18 ; give_act_reap; latency_task; check_ans;
	give_id_19 ; give_act_reap; latency_task; check_ans;
	give_id_20 ; give_act_reap; latency_task; check_ans;
	give_id_21 ; give_act_reap; latency_task; check_ans;
	give_id_22 ; give_act_reap; latency_task; check_ans;
	give_id_23 ; give_act_reap; latency_task; check_ans;
	give_id_24 ; give_act_reap; latency_task; check_ans;
	give_id_25 ; give_act_reap; latency_task; check_ans;
	give_id_26 ; give_act_reap; latency_task; check_ans;
	give_id_27 ; give_act_reap; latency_task; check_ans;
	give_id_28 ; give_act_reap; latency_task; check_ans;
	give_id_29 ; give_act_reap; latency_task; check_ans;
	give_id_30 ; give_act_reap; latency_task; check_ans;
	give_id_31 ; give_act_reap; latency_task; check_ans;
	give_id_32 ; give_act_reap; latency_task; check_ans;
	give_id_33 ; give_act_reap; latency_task; check_ans;
	give_id_34 ; give_act_reap; latency_task; check_ans;
	give_id_35 ; give_act_reap; latency_task; check_ans;
	give_id_36 ; give_act_reap; latency_task; check_ans;
	give_id_37 ; give_act_reap; latency_task; check_ans;
	give_id_38 ; give_act_reap; latency_task; check_ans;
	give_id_39 ; give_act_reap; latency_task; check_ans;
	give_id_40 ; give_act_reap; latency_task; check_ans;
	give_id_41 ; give_act_reap; latency_task; check_ans;
	give_id_42 ; give_act_reap; latency_task; check_ans;
	give_id_43 ; give_act_reap; latency_task; check_ans;
	give_id_44 ; give_act_reap; latency_task; check_ans;
	give_id_45 ; give_act_reap; latency_task; check_ans;
	give_id_46 ; give_act_reap; latency_task; check_ans;
	give_id_47 ; give_act_reap; latency_task; check_ans;
	give_id_48 ; give_act_reap; latency_task; check_ans;
	give_id_49 ; give_act_reap; latency_task; check_ans;
	give_id_50 ; give_act_reap; latency_task; check_ans;
	give_id_51 ; give_act_reap; latency_task; check_ans;
	give_id_52 ; give_act_reap; latency_task; check_ans;
	give_id_53 ; give_act_reap; latency_task; check_ans;
	give_id_54 ; give_act_reap; latency_task; check_ans;
	give_id_55 ; give_act_reap; latency_task; check_ans;
	give_id_56 ; give_act_reap; latency_task; check_ans;
	give_id_57 ; give_act_reap; latency_task; check_ans;
	give_id_58 ; give_act_reap; latency_task; check_ans;
	give_id_59 ; give_act_reap; latency_task; check_ans;
	give_id_60 ; give_act_reap; latency_task; check_ans;
	give_id_61 ; give_act_reap; latency_task; check_ans;
	give_id_62 ; give_act_reap; latency_task; check_ans;
	give_id_63 ; give_act_reap; latency_task; check_ans;
	give_id_64 ; give_act_reap; latency_task; check_ans;
	give_id_65 ; give_act_reap; latency_task; check_ans;
	give_id_66 ; give_act_reap; latency_task; check_ans;
	give_id_67 ; give_act_reap; latency_task; check_ans;
	give_id_68 ; give_act_reap; latency_task; check_ans;
	give_id_69 ; give_act_reap; latency_task; check_ans;
	give_id_70 ; give_act_reap; latency_task; check_ans;
	give_id_71 ; give_act_reap; latency_task; check_ans;
	give_id_72 ; give_act_reap; latency_task; check_ans;
	give_id_73 ; give_act_reap; latency_task; check_ans;
	give_id_74 ; give_act_reap; latency_task; check_ans;
	give_id_75 ; give_act_reap; latency_task; check_ans;
	give_id_76 ; give_act_reap; latency_task; check_ans;
	give_id_77 ; give_act_reap; latency_task; check_ans;
	give_id_78 ; give_act_reap; latency_task; check_ans;
	give_id_79 ; give_act_reap; latency_task; check_ans;
	give_id_80 ; give_act_reap; latency_task; check_ans;
	give_id_81 ; give_act_reap; latency_task; check_ans;
	give_id_82 ; give_act_reap; latency_task; check_ans;
	give_id_83 ; give_act_reap; latency_task; check_ans;
	give_id_84 ; give_act_reap; latency_task; check_ans;
	give_id_85 ; give_act_reap; latency_task; check_ans;
	give_id_86 ; give_act_reap; latency_task; check_ans;
	give_id_87 ; give_act_reap; latency_task; check_ans;
	give_id_88 ; give_act_reap; latency_task; check_ans;
	give_id_89 ; give_act_reap; latency_task; check_ans;
	give_id_90 ; give_act_reap; latency_task; check_ans;
	give_id_91 ; give_act_reap; latency_task; check_ans;
	give_id_92 ; give_act_reap; latency_task; check_ans;
	give_id_93 ; give_act_reap; latency_task; check_ans;
	give_id_94 ; give_act_reap; latency_task; check_ans;
	give_id_95 ; give_act_reap; latency_task; check_ans;
	give_id_96 ; give_act_reap; latency_task; check_ans;
	give_id_97 ; give_act_reap; latency_task; check_ans;
	give_id_98 ; give_act_reap; latency_task; check_ans;
	give_id_99 ; give_act_reap; latency_task; check_ans;
	give_id_100; give_act_reap; latency_task; check_ans;
	give_id_101; give_act_reap; latency_task; check_ans;
	give_id_102; give_act_reap; latency_task; check_ans;
	give_id_103; give_act_reap; latency_task; check_ans;
	give_id_104; give_act_reap; latency_task; check_ans;
	give_id_105; give_act_reap; latency_task; check_ans;
	give_id_106; give_act_reap; latency_task; check_ans;
	give_id_107; give_act_reap; latency_task; check_ans;
	give_id_108; give_act_reap; latency_task; check_ans;
	give_id_109; give_act_reap; latency_task; check_ans;
	give_id_110; give_act_reap; latency_task; check_ans;
	give_id_111; give_act_reap; latency_task; check_ans;
	give_id_112; give_act_reap; latency_task; check_ans;
	give_id_113; give_act_reap; latency_task; check_ans;
	give_id_114; give_act_reap; latency_task; check_ans;
	give_id_115; give_act_reap; latency_task; check_ans;
	give_id_116; give_act_reap; latency_task; check_ans;
	give_id_117; give_act_reap; latency_task; check_ans;
	give_id_118; give_act_reap; latency_task; check_ans;
	give_id_119; give_act_reap; latency_task; check_ans;
	give_id_120; give_act_reap; latency_task; check_ans;
	give_id_121; give_act_reap; latency_task; check_ans;
	give_id_122; give_act_reap; latency_task; check_ans;
	give_id_123; give_act_reap; latency_task; check_ans;
	give_id_124; give_act_reap; latency_task; check_ans;
	give_id_125; give_act_reap; latency_task; check_ans;
	give_id_126; give_act_reap; latency_task; check_ans;
	give_id_127; give_act_reap; latency_task; check_ans;
	give_id_128; give_act_reap; latency_task; check_ans;
	give_id_129; give_act_reap; latency_task; check_ans;
	give_id_130; give_act_reap; latency_task; check_ans;
	give_id_131; give_act_reap; latency_task; check_ans;
	give_id_132; give_act_reap; latency_task; check_ans;
	give_id_133; give_act_reap; latency_task; check_ans;
	give_id_134; give_act_reap; latency_task; check_ans;
	give_id_135; give_act_reap; latency_task; check_ans;
	give_id_136; give_act_reap; latency_task; check_ans;
	give_id_137; give_act_reap; latency_task; check_ans;
	give_id_138; give_act_reap; latency_task; check_ans;
	give_id_139; give_act_reap; latency_task; check_ans;
	give_id_140; give_act_reap; latency_task; check_ans;
	give_id_141; give_act_reap; latency_task; check_ans;
	give_id_142; give_act_reap; latency_task; check_ans;
	give_id_143; give_act_reap; latency_task; check_ans;
	give_id_144; give_act_reap; latency_task; check_ans;
	give_id_145; give_act_reap; latency_task; check_ans;
	give_id_146; give_act_reap; latency_task; check_ans;
	give_id_147; give_act_reap; latency_task; check_ans;
	give_id_148; give_act_reap; latency_task; check_ans;
	give_id_149; give_act_reap; latency_task; check_ans;
	give_id_150; give_act_reap; latency_task; check_ans;
	give_id_151; give_act_reap; latency_task; check_ans;
	give_id_152; give_act_reap; latency_task; check_ans;
	give_id_153; give_act_reap; latency_task; check_ans;
	give_id_154; give_act_reap; latency_task; check_ans;
	give_id_155; give_act_reap; latency_task; check_ans;
	give_id_156; give_act_reap; latency_task; check_ans;
	give_id_157; give_act_reap; latency_task; check_ans;
	give_id_158; give_act_reap; latency_task; check_ans;
	give_id_159; give_act_reap; latency_task; check_ans;
	give_id_160; give_act_reap; latency_task; check_ans;
	give_id_161; give_act_reap; latency_task; check_ans;
	give_id_162; give_act_reap; latency_task; check_ans;
	give_id_163; give_act_reap; latency_task; check_ans;
	give_id_164; give_act_reap; latency_task; check_ans;
	give_id_165; give_act_reap; latency_task; check_ans;
	give_id_166; give_act_reap; latency_task; check_ans;
	give_id_167; give_act_reap; latency_task; check_ans;
	give_id_168; give_act_reap; latency_task; check_ans;
	give_id_169; give_act_reap; latency_task; check_ans;
	give_id_170; give_act_reap; latency_task; check_ans;
	give_id_171; give_act_reap; latency_task; check_ans;
	give_id_172; give_act_reap; latency_task; check_ans;
	give_id_173; give_act_reap; latency_task; check_ans;
	give_id_174; give_act_reap; latency_task; check_ans;
	give_id_175; give_act_reap; latency_task; check_ans;
	give_id_176; give_act_reap; latency_task; check_ans;
	give_id_177; give_act_reap; latency_task; check_ans;
	give_id_178; give_act_reap; latency_task; check_ans;
	give_id_179; give_act_reap; latency_task; check_ans;
	give_id_180; give_act_reap; latency_task; check_ans;
	give_id_181; give_act_reap; latency_task; check_ans;
	give_id_182; give_act_reap; latency_task; check_ans;
	give_id_183; give_act_reap; latency_task; check_ans;
	give_id_184; give_act_reap; latency_task; check_ans;
	give_id_185; give_act_reap; latency_task; check_ans;
	give_id_186; give_act_reap; latency_task; check_ans;
	give_id_187; give_act_reap; latency_task; check_ans;
	give_id_188; give_act_reap; latency_task; check_ans;
	give_id_189; give_act_reap; latency_task; check_ans;
	give_id_190; give_act_reap; latency_task; check_ans;
	give_id_191; give_act_reap; latency_task; check_ans;
	give_id_192; give_act_reap; latency_task; check_ans;
	give_id_193; give_act_reap; latency_task; check_ans;
	give_id_194; give_act_reap; latency_task; check_ans;
	give_id_195; give_act_reap; latency_task; check_ans;
	give_id_196; give_act_reap; latency_task; check_ans;
	give_id_197; give_act_reap; latency_task; check_ans;
	give_id_198; give_act_reap; latency_task; check_ans;
	give_id_199; give_act_reap; latency_task; check_ans;
	give_id_200; give_act_reap; latency_task; check_ans;
	give_id_201; give_act_reap; latency_task; check_ans;
	give_id_202; give_act_reap; latency_task; check_ans;
	give_id_203; give_act_reap; latency_task; check_ans;
	give_id_204; give_act_reap; latency_task; check_ans;
	give_id_205; give_act_reap; latency_task; check_ans;
	give_id_206; give_act_reap; latency_task; check_ans;
	give_id_207; give_act_reap; latency_task; check_ans;
	give_id_208; give_act_reap; latency_task; check_ans;
	give_id_209; give_act_reap; latency_task; check_ans;
	give_id_210; give_act_reap; latency_task; check_ans;
	give_id_211; give_act_reap; latency_task; check_ans;
	give_id_212; give_act_reap; latency_task; check_ans;
	give_id_213; give_act_reap; latency_task; check_ans;
	give_id_214; give_act_reap; latency_task; check_ans;
	give_id_215; give_act_reap; latency_task; check_ans;
	give_id_216; give_act_reap; latency_task; check_ans;
	give_id_217; give_act_reap; latency_task; check_ans;
	give_id_218; give_act_reap; latency_task; check_ans;
	give_id_219; give_act_reap; latency_task; check_ans;
	give_id_220; give_act_reap; latency_task; check_ans;
	give_id_221; give_act_reap; latency_task; check_ans;
	give_id_222; give_act_reap; latency_task; check_ans;
	give_id_223; give_act_reap; latency_task; check_ans;
	give_id_224; give_act_reap; latency_task; check_ans;
	give_id_225; give_act_reap; latency_task; check_ans;
	give_id_226; give_act_reap; latency_task; check_ans;
	give_id_227; give_act_reap; latency_task; check_ans;
	give_id_228; give_act_reap; latency_task; check_ans;
	give_id_229; give_act_reap; latency_task; check_ans;
	give_id_230; give_act_reap; latency_task; check_ans;
	give_id_231; give_act_reap; latency_task; check_ans;
	give_id_232; give_act_reap; latency_task; check_ans;
	give_id_233; give_act_reap; latency_task; check_ans;
	give_id_234; give_act_reap; latency_task; check_ans;
	give_id_235; give_act_reap; latency_task; check_ans;
	give_id_236; give_act_reap; latency_task; check_ans;
	give_id_237; give_act_reap; latency_task; check_ans;
	give_id_238; give_act_reap; latency_task; check_ans;
	give_id_239; give_act_reap; latency_task; check_ans;
	give_id_240; give_act_reap; latency_task; check_ans;
	give_id_241; give_act_reap; latency_task; check_ans;
	give_id_242; give_act_reap; latency_task; check_ans;
	give_id_243; give_act_reap; latency_task; check_ans;
	give_id_244; give_act_reap; latency_task; check_ans;
	give_id_245; give_act_reap; latency_task; check_ans;
	give_id_246; give_act_reap; latency_task; check_ans;
	give_id_247; give_act_reap; latency_task; check_ans;
	give_id_248; give_act_reap; latency_task; check_ans;
	give_id_249; give_act_reap; latency_task; check_ans;
	give_id_250; give_act_reap; latency_task; check_ans;
	give_id_251; give_act_reap; latency_task; check_ans;
	give_id_252; give_act_reap; latency_task; check_ans;
	give_id_253; give_act_reap; latency_task; check_ans;
	give_id_254; give_act_reap; latency_task; check_ans;
	// ID 9
	give_id_0  ; give_act_reap; latency_task; check_ans;
	give_id_1  ; give_act_reap; latency_task; check_ans;
	give_id_2  ; give_act_reap; latency_task; check_ans;
	give_id_3  ; give_act_reap; latency_task; check_ans;
	give_id_4  ; give_act_reap; latency_task; check_ans;
	give_id_5  ; give_act_reap; latency_task; check_ans;
	give_id_6  ; give_act_reap; latency_task; check_ans;
	give_id_7  ; give_act_reap; latency_task; check_ans;
	give_id_8  ; give_act_reap; latency_task; check_ans;
	give_id_9  ; give_act_reap; latency_task; check_ans;
	give_id_10 ; give_act_reap; latency_task; check_ans;
	give_id_11 ; give_act_reap; latency_task; check_ans;
	give_id_12 ; give_act_reap; latency_task; check_ans;
	give_id_13 ; give_act_reap; latency_task; check_ans;
	give_id_14 ; give_act_reap; latency_task; check_ans;
	give_id_15 ; give_act_reap; latency_task; check_ans;
	give_id_16 ; give_act_reap; latency_task; check_ans;
	give_id_17 ; give_act_reap; latency_task; check_ans;
	give_id_18 ; give_act_reap; latency_task; check_ans;
	give_id_19 ; give_act_reap; latency_task; check_ans;
	give_id_20 ; give_act_reap; latency_task; check_ans;
	give_id_21 ; give_act_reap; latency_task; check_ans;
	give_id_22 ; give_act_reap; latency_task; check_ans;
	give_id_23 ; give_act_reap; latency_task; check_ans;
	give_id_24 ; give_act_reap; latency_task; check_ans;
	give_id_25 ; give_act_reap; latency_task; check_ans;
	give_id_26 ; give_act_reap; latency_task; check_ans;
	give_id_27 ; give_act_reap; latency_task; check_ans;
	give_id_28 ; give_act_reap; latency_task; check_ans;
	give_id_29 ; give_act_reap; latency_task; check_ans;
	give_id_30 ; give_act_reap; latency_task; check_ans;
	give_id_31 ; give_act_reap; latency_task; check_ans;
	give_id_32 ; give_act_reap; latency_task; check_ans;
	give_id_33 ; give_act_reap; latency_task; check_ans;
	give_id_34 ; give_act_reap; latency_task; check_ans;
	give_id_35 ; give_act_reap; latency_task; check_ans;
	give_id_36 ; give_act_reap; latency_task; check_ans;
	give_id_37 ; give_act_reap; latency_task; check_ans;
	give_id_38 ; give_act_reap; latency_task; check_ans;
	give_id_39 ; give_act_reap; latency_task; check_ans;
	give_id_40 ; give_act_reap; latency_task; check_ans;
	give_id_41 ; give_act_reap; latency_task; check_ans;
	give_id_42 ; give_act_reap; latency_task; check_ans;
	give_id_43 ; give_act_reap; latency_task; check_ans;
	give_id_44 ; give_act_reap; latency_task; check_ans;
	give_id_45 ; give_act_reap; latency_task; check_ans;
	give_id_46 ; give_act_reap; latency_task; check_ans;
	give_id_47 ; give_act_reap; latency_task; check_ans;
	give_id_48 ; give_act_reap; latency_task; check_ans;
	give_id_49 ; give_act_reap; latency_task; check_ans;
	give_id_50 ; give_act_reap; latency_task; check_ans;
	give_id_51 ; give_act_reap; latency_task; check_ans;
	give_id_52 ; give_act_reap; latency_task; check_ans;
	give_id_53 ; give_act_reap; latency_task; check_ans;
	give_id_54 ; give_act_reap; latency_task; check_ans;
	give_id_55 ; give_act_reap; latency_task; check_ans;
	give_id_56 ; give_act_reap; latency_task; check_ans;
	give_id_57 ; give_act_reap; latency_task; check_ans;
	give_id_58 ; give_act_reap; latency_task; check_ans;
	give_id_59 ; give_act_reap; latency_task; check_ans;
	give_id_60 ; give_act_reap; latency_task; check_ans;
	give_id_61 ; give_act_reap; latency_task; check_ans;
	give_id_62 ; give_act_reap; latency_task; check_ans;
	give_id_63 ; give_act_reap; latency_task; check_ans;
	give_id_64 ; give_act_reap; latency_task; check_ans;
	give_id_65 ; give_act_reap; latency_task; check_ans;
	give_id_66 ; give_act_reap; latency_task; check_ans;
	give_id_67 ; give_act_reap; latency_task; check_ans;
	give_id_68 ; give_act_reap; latency_task; check_ans;
	give_id_69 ; give_act_reap; latency_task; check_ans;
	give_id_70 ; give_act_reap; latency_task; check_ans;
	give_id_71 ; give_act_reap; latency_task; check_ans;
	give_id_72 ; give_act_reap; latency_task; check_ans;
	give_id_73 ; give_act_reap; latency_task; check_ans;
	give_id_74 ; give_act_reap; latency_task; check_ans;
	give_id_75 ; give_act_reap; latency_task; check_ans;
	give_id_76 ; give_act_reap; latency_task; check_ans;
	give_id_77 ; give_act_reap; latency_task; check_ans;
	give_id_78 ; give_act_reap; latency_task; check_ans;
	give_id_79 ; give_act_reap; latency_task; check_ans;
	give_id_80 ; give_act_reap; latency_task; check_ans;
	give_id_81 ; give_act_reap; latency_task; check_ans;
	give_id_82 ; give_act_reap; latency_task; check_ans;
	give_id_83 ; give_act_reap; latency_task; check_ans;
	give_id_84 ; give_act_reap; latency_task; check_ans;
	give_id_85 ; give_act_reap; latency_task; check_ans;
	give_id_86 ; give_act_reap; latency_task; check_ans;
	give_id_87 ; give_act_reap; latency_task; check_ans;
	give_id_88 ; give_act_reap; latency_task; check_ans;
	give_id_89 ; give_act_reap; latency_task; check_ans;
	give_id_90 ; give_act_reap; latency_task; check_ans;
	give_id_91 ; give_act_reap; latency_task; check_ans;
	give_id_92 ; give_act_reap; latency_task; check_ans;
	give_id_93 ; give_act_reap; latency_task; check_ans;
	give_id_94 ; give_act_reap; latency_task; check_ans;
	give_id_95 ; give_act_reap; latency_task; check_ans;
	give_id_96 ; give_act_reap; latency_task; check_ans;
	give_id_97 ; give_act_reap; latency_task; check_ans;
	give_id_98 ; give_act_reap; latency_task; check_ans;
	give_id_99 ; give_act_reap; latency_task; check_ans;
	give_id_100; give_act_reap; latency_task; check_ans;
	give_id_101; give_act_reap; latency_task; check_ans;
	give_id_102; give_act_reap; latency_task; check_ans;
	give_id_103; give_act_reap; latency_task; check_ans;
	give_id_104; give_act_reap; latency_task; check_ans;
	give_id_105; give_act_reap; latency_task; check_ans;
	give_id_106; give_act_reap; latency_task; check_ans;
	give_id_107; give_act_reap; latency_task; check_ans;
	give_id_108; give_act_reap; latency_task; check_ans;
	give_id_109; give_act_reap; latency_task; check_ans;
	give_id_110; give_act_reap; latency_task; check_ans;
	give_id_111; give_act_reap; latency_task; check_ans;
	give_id_112; give_act_reap; latency_task; check_ans;
	give_id_113; give_act_reap; latency_task; check_ans;
	give_id_114; give_act_reap; latency_task; check_ans;
	give_id_115; give_act_reap; latency_task; check_ans;
	give_id_116; give_act_reap; latency_task; check_ans;
	give_id_117; give_act_reap; latency_task; check_ans;
	give_id_118; give_act_reap; latency_task; check_ans;
	give_id_119; give_act_reap; latency_task; check_ans;
	give_id_120; give_act_reap; latency_task; check_ans;
	give_id_121; give_act_reap; latency_task; check_ans;
	give_id_122; give_act_reap; latency_task; check_ans;
	give_id_123; give_act_reap; latency_task; check_ans;
	give_id_124; give_act_reap; latency_task; check_ans;
	give_id_125; give_act_reap; latency_task; check_ans;
	give_id_126; give_act_reap; latency_task; check_ans;
	give_id_127; give_act_reap; latency_task; check_ans;
	give_id_128; give_act_reap; latency_task; check_ans;
	give_id_129; give_act_reap; latency_task; check_ans;
	give_id_130; give_act_reap; latency_task; check_ans;
	give_id_131; give_act_reap; latency_task; check_ans;
	give_id_132; give_act_reap; latency_task; check_ans;
	give_id_133; give_act_reap; latency_task; check_ans;
	give_id_134; give_act_reap; latency_task; check_ans;
	give_id_135; give_act_reap; latency_task; check_ans;
	give_id_136; give_act_reap; latency_task; check_ans;
	give_id_137; give_act_reap; latency_task; check_ans;
	give_id_138; give_act_reap; latency_task; check_ans;
	give_id_139; give_act_reap; latency_task; check_ans;
	give_id_140; give_act_reap; latency_task; check_ans;
	give_id_141; give_act_reap; latency_task; check_ans;
	give_id_142; give_act_reap; latency_task; check_ans;
	give_id_143; give_act_reap; latency_task; check_ans;
	give_id_144; give_act_reap; latency_task; check_ans;
	give_id_145; give_act_reap; latency_task; check_ans;
	give_id_146; give_act_reap; latency_task; check_ans;
	give_id_147; give_act_reap; latency_task; check_ans;
	give_id_148; give_act_reap; latency_task; check_ans;
	give_id_149; give_act_reap; latency_task; check_ans;
	give_id_150; give_act_reap; latency_task; check_ans;
	give_id_151; give_act_reap; latency_task; check_ans;
	give_id_152; give_act_reap; latency_task; check_ans;
	give_id_153; give_act_reap; latency_task; check_ans;
	give_id_154; give_act_reap; latency_task; check_ans;
	give_id_155; give_act_reap; latency_task; check_ans;
	give_id_156; give_act_reap; latency_task; check_ans;
	give_id_157; give_act_reap; latency_task; check_ans;
	give_id_158; give_act_reap; latency_task; check_ans;
	give_id_159; give_act_reap; latency_task; check_ans;
	give_id_160; give_act_reap; latency_task; check_ans;
	give_id_161; give_act_reap; latency_task; check_ans;
	give_id_162; give_act_reap; latency_task; check_ans;
	give_id_163; give_act_reap; latency_task; check_ans;
	give_id_164; give_act_reap; latency_task; check_ans;
	give_id_165; give_act_reap; latency_task; check_ans;
	give_id_166; give_act_reap; latency_task; check_ans;
	give_id_167; give_act_reap; latency_task; check_ans;
	give_id_168; give_act_reap; latency_task; check_ans;
	give_id_169; give_act_reap; latency_task; check_ans;
	give_id_170; give_act_reap; latency_task; check_ans;
	give_id_171; give_act_reap; latency_task; check_ans;
	give_id_172; give_act_reap; latency_task; check_ans;
	give_id_173; give_act_reap; latency_task; check_ans;
	give_id_174; give_act_reap; latency_task; check_ans;
	give_id_175; give_act_reap; latency_task; check_ans;
	give_id_176; give_act_reap; latency_task; check_ans;
	give_id_177; give_act_reap; latency_task; check_ans;
	give_id_178; give_act_reap; latency_task; check_ans;
	give_id_179; give_act_reap; latency_task; check_ans;
	give_id_180; give_act_reap; latency_task; check_ans;
	give_id_181; give_act_reap; latency_task; check_ans;
	give_id_182; give_act_reap; latency_task; check_ans;
	give_id_183; give_act_reap; latency_task; check_ans;
	give_id_184; give_act_reap; latency_task; check_ans;
	give_id_185; give_act_reap; latency_task; check_ans;
	give_id_186; give_act_reap; latency_task; check_ans;
	give_id_187; give_act_reap; latency_task; check_ans;
	give_id_188; give_act_reap; latency_task; check_ans;
	give_id_189; give_act_reap; latency_task; check_ans;
	give_id_190; give_act_reap; latency_task; check_ans;
	give_id_191; give_act_reap; latency_task; check_ans;
	give_id_192; give_act_reap; latency_task; check_ans;
	give_id_193; give_act_reap; latency_task; check_ans;
	give_id_194; give_act_reap; latency_task; check_ans;
	give_id_195; give_act_reap; latency_task; check_ans;
	give_id_196; give_act_reap; latency_task; check_ans;
	give_id_197; give_act_reap; latency_task; check_ans;
	give_id_198; give_act_reap; latency_task; check_ans;
	give_id_199; give_act_reap; latency_task; check_ans;
	give_id_200; give_act_reap; latency_task; check_ans;
	give_id_201; give_act_reap; latency_task; check_ans;
	give_id_202; give_act_reap; latency_task; check_ans;
	give_id_203; give_act_reap; latency_task; check_ans;
	give_id_204; give_act_reap; latency_task; check_ans;
	give_id_205; give_act_reap; latency_task; check_ans;
	give_id_206; give_act_reap; latency_task; check_ans;
	give_id_207; give_act_reap; latency_task; check_ans;
	give_id_208; give_act_reap; latency_task; check_ans;
	give_id_209; give_act_reap; latency_task; check_ans;
	give_id_210; give_act_reap; latency_task; check_ans;
	give_id_211; give_act_reap; latency_task; check_ans;
	give_id_212; give_act_reap; latency_task; check_ans;
	give_id_213; give_act_reap; latency_task; check_ans;
	give_id_214; give_act_reap; latency_task; check_ans;
	give_id_215; give_act_reap; latency_task; check_ans;
	give_id_216; give_act_reap; latency_task; check_ans;
	give_id_217; give_act_reap; latency_task; check_ans;
	give_id_218; give_act_reap; latency_task; check_ans;
	give_id_219; give_act_reap; latency_task; check_ans;
	give_id_220; give_act_reap; latency_task; check_ans;
	give_id_221; give_act_reap; latency_task; check_ans;
	give_id_222; give_act_reap; latency_task; check_ans;
	give_id_223; give_act_reap; latency_task; check_ans;
	give_id_224; give_act_reap; latency_task; check_ans;
	give_id_225; give_act_reap; latency_task; check_ans;
	give_id_226; give_act_reap; latency_task; check_ans;
	give_id_227; give_act_reap; latency_task; check_ans;
	give_id_228; give_act_reap; latency_task; check_ans;
	give_id_229; give_act_reap; latency_task; check_ans;
	give_id_230; give_act_reap; latency_task; check_ans;
	give_id_231; give_act_reap; latency_task; check_ans;
	give_id_232; give_act_reap; latency_task; check_ans;
	give_id_233; give_act_reap; latency_task; check_ans;
	give_id_234; give_act_reap; latency_task; check_ans;
	give_id_235; give_act_reap; latency_task; check_ans;
	give_id_236; give_act_reap; latency_task; check_ans;
	give_id_237; give_act_reap; latency_task; check_ans;
	give_id_238; give_act_reap; latency_task; check_ans;
	give_id_239; give_act_reap; latency_task; check_ans;
	give_id_240; give_act_reap; latency_task; check_ans;
	give_id_241; give_act_reap; latency_task; check_ans;
	give_id_242; give_act_reap; latency_task; check_ans;
	give_id_243; give_act_reap; latency_task; check_ans;
	give_id_244; give_act_reap; latency_task; check_ans;
	give_id_245; give_act_reap; latency_task; check_ans;
	give_id_246; give_act_reap; latency_task; check_ans;
	give_id_247; give_act_reap; latency_task; check_ans;
	give_id_248; give_act_reap; latency_task; check_ans;
	give_id_249; give_act_reap; latency_task; check_ans;
	give_id_250; give_act_reap; latency_task; check_ans;
	give_id_251; give_act_reap; latency_task; check_ans;
	give_id_252; give_act_reap; latency_task; check_ans;
	give_id_253; give_act_reap; latency_task; check_ans;
	give_id_254; give_act_reap; latency_task; check_ans;
	// ID 10
	give_id_0  ; give_act_reap; latency_task; check_ans;
	give_id_1  ; give_act_reap; latency_task; check_ans;
	give_id_2  ; give_act_reap; latency_task; check_ans;
	give_id_3  ; give_act_reap; latency_task; check_ans;
	give_id_4  ; give_act_reap; latency_task; check_ans;
	give_id_5  ; give_act_reap; latency_task; check_ans;
	give_id_6  ; give_act_reap; latency_task; check_ans;
	give_id_7  ; give_act_reap; latency_task; check_ans;
	give_id_8  ; give_act_reap; latency_task; check_ans;
	give_id_9  ; give_act_reap; latency_task; check_ans;
	give_id_10 ; give_act_reap; latency_task; check_ans;
	give_id_11 ; give_act_reap; latency_task; check_ans;
	give_id_12 ; give_act_reap; latency_task; check_ans;
	give_id_13 ; give_act_reap; latency_task; check_ans;
	give_id_14 ; give_act_reap; latency_task; check_ans;
	give_id_15 ; give_act_reap; latency_task; check_ans;
	give_id_16 ; give_act_reap; latency_task; check_ans;
	give_id_17 ; give_act_reap; latency_task; check_ans;
	give_id_18 ; give_act_reap; latency_task; check_ans;
	give_id_19 ; give_act_reap; latency_task; check_ans;
	give_id_20 ; give_act_reap; latency_task; check_ans;
	give_id_21 ; give_act_reap; latency_task; check_ans;
	give_id_22 ; give_act_reap; latency_task; check_ans;
	give_id_23 ; give_act_reap; latency_task; check_ans;
	give_id_24 ; give_act_reap; latency_task; check_ans;
	give_id_25 ; give_act_reap; latency_task; check_ans;
	give_id_26 ; give_act_reap; latency_task; check_ans;
	give_id_27 ; give_act_reap; latency_task; check_ans;
	give_id_28 ; give_act_reap; latency_task; check_ans;
	give_id_29 ; give_act_reap; latency_task; check_ans;
	give_id_30 ; give_act_reap; latency_task; check_ans;
	give_id_31 ; give_act_reap; latency_task; check_ans;
	give_id_32 ; give_act_reap; latency_task; check_ans;
	give_id_33 ; give_act_reap; latency_task; check_ans;
	give_id_34 ; give_act_reap; latency_task; check_ans;
	give_id_35 ; give_act_reap; latency_task; check_ans;
	give_id_36 ; give_act_reap; latency_task; check_ans;
	give_id_37 ; give_act_reap; latency_task; check_ans;
	give_id_38 ; give_act_reap; latency_task; check_ans;
	give_id_39 ; give_act_reap; latency_task; check_ans;
	give_id_40 ; give_act_reap; latency_task; check_ans;
	give_id_41 ; give_act_reap; latency_task; check_ans;
	give_id_42 ; give_act_reap; latency_task; check_ans;
	give_id_43 ; give_act_reap; latency_task; check_ans;
	give_id_44 ; give_act_reap; latency_task; check_ans;
	give_id_45 ; give_act_reap; latency_task; check_ans;
	give_id_46 ; give_act_reap; latency_task; check_ans;
	give_id_47 ; give_act_reap; latency_task; check_ans;
	give_id_48 ; give_act_reap; latency_task; check_ans;
	give_id_49 ; give_act_reap; latency_task; check_ans;
	give_id_50 ; give_act_reap; latency_task; check_ans;
	give_id_51 ; give_act_reap; latency_task; check_ans;
	give_id_52 ; give_act_reap; latency_task; check_ans;
	give_id_53 ; give_act_reap; latency_task; check_ans;
	give_id_54 ; give_act_reap; latency_task; check_ans;
	give_id_55 ; give_act_reap; latency_task; check_ans;
	give_id_56 ; give_act_reap; latency_task; check_ans;
	give_id_57 ; give_act_reap; latency_task; check_ans;
	give_id_58 ; give_act_reap; latency_task; check_ans;
	give_id_59 ; give_act_reap; latency_task; check_ans;
	give_id_60 ; give_act_reap; latency_task; check_ans;
	give_id_61 ; give_act_reap; latency_task; check_ans;
	give_id_62 ; give_act_reap; latency_task; check_ans;
	give_id_63 ; give_act_reap; latency_task; check_ans;
	give_id_64 ; give_act_reap; latency_task; check_ans;
	give_id_65 ; give_act_reap; latency_task; check_ans;
	give_id_66 ; give_act_reap; latency_task; check_ans;
	give_id_67 ; give_act_reap; latency_task; check_ans;
	give_id_68 ; give_act_reap; latency_task; check_ans;
	give_id_69 ; give_act_reap; latency_task; check_ans;
	give_id_70 ; give_act_reap; latency_task; check_ans;
	give_id_71 ; give_act_reap; latency_task; check_ans;
	give_id_72 ; give_act_reap; latency_task; check_ans;
	give_id_73 ; give_act_reap; latency_task; check_ans;
	give_id_74 ; give_act_reap; latency_task; check_ans;
	give_id_75 ; give_act_reap; latency_task; check_ans;
	give_id_76 ; give_act_reap; latency_task; check_ans;
	give_id_77 ; give_act_reap; latency_task; check_ans;
	give_id_78 ; give_act_reap; latency_task; check_ans;
	give_id_79 ; give_act_reap; latency_task; check_ans;
	give_id_80 ; give_act_reap; latency_task; check_ans;
	give_id_81 ; give_act_reap; latency_task; check_ans;
	give_id_82 ; give_act_reap; latency_task; check_ans;
	give_id_83 ; give_act_reap; latency_task; check_ans;
	give_id_84 ; give_act_reap; latency_task; check_ans;
	give_id_85 ; give_act_reap; latency_task; check_ans;
	give_id_86 ; give_act_reap; latency_task; check_ans;
	give_id_87 ; give_act_reap; latency_task; check_ans;
	give_id_88 ; give_act_reap; latency_task; check_ans;
	give_id_89 ; give_act_reap; latency_task; check_ans;
	give_id_90 ; give_act_reap; latency_task; check_ans;
	give_id_91 ; give_act_reap; latency_task; check_ans;
	give_id_92 ; give_act_reap; latency_task; check_ans;
	give_id_93 ; give_act_reap; latency_task; check_ans;
	give_id_94 ; give_act_reap; latency_task; check_ans;
	give_id_95 ; give_act_reap; latency_task; check_ans;
	give_id_96 ; give_act_reap; latency_task; check_ans;
	give_id_97 ; give_act_reap; latency_task; check_ans;
	give_id_98 ; give_act_reap; latency_task; check_ans;
	give_id_99 ; give_act_reap; latency_task; check_ans;
	give_id_100; give_act_reap; latency_task; check_ans;
	give_id_101; give_act_reap; latency_task; check_ans;
	give_id_102; give_act_reap; latency_task; check_ans;
	give_id_103; give_act_reap; latency_task; check_ans;
	give_id_104; give_act_reap; latency_task; check_ans;
	give_id_105; give_act_reap; latency_task; check_ans;
	give_id_106; give_act_reap; latency_task; check_ans;
	give_id_107; give_act_reap; latency_task; check_ans;
	give_id_108; give_act_reap; latency_task; check_ans;
	give_id_109; give_act_reap; latency_task; check_ans;
	give_id_110; give_act_reap; latency_task; check_ans;
	give_id_111; give_act_reap; latency_task; check_ans;
	give_id_112; give_act_reap; latency_task; check_ans;
	give_id_113; give_act_reap; latency_task; check_ans;
	give_id_114; give_act_reap; latency_task; check_ans;
	give_id_115; give_act_reap; latency_task; check_ans;
	give_id_116; give_act_reap; latency_task; check_ans;
	give_id_117; give_act_reap; latency_task; check_ans;
	give_id_118; give_act_reap; latency_task; check_ans;
	give_id_119; give_act_reap; latency_task; check_ans;
	give_id_120; give_act_reap; latency_task; check_ans;
	give_id_121; give_act_reap; latency_task; check_ans;
	give_id_122; give_act_reap; latency_task; check_ans;
	give_id_123; give_act_reap; latency_task; check_ans;
	give_id_124; give_act_reap; latency_task; check_ans;
	give_id_125; give_act_reap; latency_task; check_ans;
	give_id_126; give_act_reap; latency_task; check_ans;
	give_id_127; give_act_reap; latency_task; check_ans;
	give_id_128; give_act_reap; latency_task; check_ans;
	give_id_129; give_act_reap; latency_task; check_ans;
	give_id_130; give_act_reap; latency_task; check_ans;
	give_id_131; give_act_reap; latency_task; check_ans;
	give_id_132; give_act_reap; latency_task; check_ans;
	give_id_133; give_act_reap; latency_task; check_ans;
	give_id_134; give_act_reap; latency_task; check_ans;
	give_id_135; give_act_reap; latency_task; check_ans;
	give_id_136; give_act_reap; latency_task; check_ans;
	give_id_137; give_act_reap; latency_task; check_ans;
	give_id_138; give_act_reap; latency_task; check_ans;
	give_id_139; give_act_reap; latency_task; check_ans;
	give_id_140; give_act_reap; latency_task; check_ans;
	give_id_141; give_act_reap; latency_task; check_ans;
	give_id_142; give_act_reap; latency_task; check_ans;
	give_id_143; give_act_reap; latency_task; check_ans;
	give_id_144; give_act_reap; latency_task; check_ans;
	give_id_145; give_act_reap; latency_task; check_ans;
	give_id_146; give_act_reap; latency_task; check_ans;
	give_id_147; give_act_reap; latency_task; check_ans;
	give_id_148; give_act_reap; latency_task; check_ans;
	give_id_149; give_act_reap; latency_task; check_ans;
	give_id_150; give_act_reap; latency_task; check_ans;
	give_id_151; give_act_reap; latency_task; check_ans;
	give_id_152; give_act_reap; latency_task; check_ans;
	give_id_153; give_act_reap; latency_task; check_ans;
	give_id_154; give_act_reap; latency_task; check_ans;
	give_id_155; give_act_reap; latency_task; check_ans;
	give_id_156; give_act_reap; latency_task; check_ans;
	give_id_157; give_act_reap; latency_task; check_ans;
	give_id_158; give_act_reap; latency_task; check_ans;
	give_id_159; give_act_reap; latency_task; check_ans;
	give_id_160; give_act_reap; latency_task; check_ans;
	give_id_161; give_act_reap; latency_task; check_ans;
	give_id_162; give_act_reap; latency_task; check_ans;
	give_id_163; give_act_reap; latency_task; check_ans;
	give_id_164; give_act_reap; latency_task; check_ans;
	give_id_165; give_act_reap; latency_task; check_ans;
	give_id_166; give_act_reap; latency_task; check_ans;
	give_id_167; give_act_reap; latency_task; check_ans;
	give_id_168; give_act_reap; latency_task; check_ans;
	give_id_169; give_act_reap; latency_task; check_ans;
	give_id_170; give_act_reap; latency_task; check_ans;
	give_id_171; give_act_reap; latency_task; check_ans;
	give_id_172; give_act_reap; latency_task; check_ans;
	give_id_173; give_act_reap; latency_task; check_ans;
	give_id_174; give_act_reap; latency_task; check_ans;
	give_id_175; give_act_reap; latency_task; check_ans;
	give_id_176; give_act_reap; latency_task; check_ans;
	give_id_177; give_act_reap; latency_task; check_ans;
	give_id_178; give_act_reap; latency_task; check_ans;
	give_id_179; give_act_reap; latency_task; check_ans;
	give_id_180; give_act_reap; latency_task; check_ans;
	give_id_181; give_act_reap; latency_task; check_ans;
	give_id_182; give_act_reap; latency_task; check_ans;
	give_id_183; give_act_reap; latency_task; check_ans;
	give_id_184; give_act_reap; latency_task; check_ans;
	give_id_185; give_act_reap; latency_task; check_ans;
	give_id_186; give_act_reap; latency_task; check_ans;
	give_id_187; give_act_reap; latency_task; check_ans;
	give_id_188; give_act_reap; latency_task; check_ans;
	give_id_189; give_act_reap; latency_task; check_ans;
	give_id_190; give_act_reap; latency_task; check_ans;
	give_id_191; give_act_reap; latency_task; check_ans;
	give_id_192; give_act_reap; latency_task; check_ans;
	give_id_193; give_act_reap; latency_task; check_ans;
	give_id_194; give_act_reap; latency_task; check_ans;
	give_id_195; give_act_reap; latency_task; check_ans;
	give_id_196; give_act_reap; latency_task; check_ans;
	give_id_197; give_act_reap; latency_task; check_ans;
	give_id_198; give_act_reap; latency_task; check_ans;
	give_id_199; give_act_reap; latency_task; check_ans;
	give_id_200; give_act_reap; latency_task; check_ans;
	give_id_201; give_act_reap; latency_task; check_ans;
	give_id_202; give_act_reap; latency_task; check_ans;
	give_id_203; give_act_reap; latency_task; check_ans;
	give_id_204; give_act_reap; latency_task; check_ans;
	give_id_205; give_act_reap; latency_task; check_ans;
	give_id_206; give_act_reap; latency_task; check_ans;
	give_id_207; give_act_reap; latency_task; check_ans;
	give_id_208; give_act_reap; latency_task; check_ans;
	give_id_209; give_act_reap; latency_task; check_ans;
	give_id_210; give_act_reap; latency_task; check_ans;
	give_id_211; give_act_reap; latency_task; check_ans;
	give_id_212; give_act_reap; latency_task; check_ans;
	give_id_213; give_act_reap; latency_task; check_ans;
	give_id_214; give_act_reap; latency_task; check_ans;
	give_id_215; give_act_reap; latency_task; check_ans;
	give_id_216; give_act_reap; latency_task; check_ans;
	give_id_217; give_act_reap; latency_task; check_ans;
	give_id_218; give_act_reap; latency_task; check_ans;
	give_id_219; give_act_reap; latency_task; check_ans;
	give_id_220; give_act_reap; latency_task; check_ans;
	give_id_221; give_act_reap; latency_task; check_ans;
	give_id_222; give_act_reap; latency_task; check_ans;
	give_id_223; give_act_reap; latency_task; check_ans;
	give_id_224; give_act_reap; latency_task; check_ans;
	give_id_225; give_act_reap; latency_task; check_ans;
	give_id_226; give_act_reap; latency_task; check_ans;
	give_id_227; give_act_reap; latency_task; check_ans;
	give_id_228; give_act_reap; latency_task; check_ans;
	give_id_229; give_act_reap; latency_task; check_ans;
	give_id_230; give_act_reap; latency_task; check_ans;
	give_id_231; give_act_reap; latency_task; check_ans;
	give_id_232; give_act_reap; latency_task; check_ans;
	give_id_233; give_act_reap; latency_task; check_ans;
	give_id_234; give_act_reap; latency_task; check_ans;
	give_id_235; give_act_reap; latency_task; check_ans;
	give_id_236; give_act_reap; latency_task; check_ans;
	give_id_237; give_act_reap; latency_task; check_ans;
	give_id_238; give_act_reap; latency_task; check_ans;
	give_id_239; give_act_reap; latency_task; check_ans;
	give_id_240; give_act_reap; latency_task; check_ans;
	give_id_241; give_act_reap; latency_task; check_ans;
	give_id_242; give_act_reap; latency_task; check_ans;
	give_id_243; give_act_reap; latency_task; check_ans;
	give_id_244; give_act_reap; latency_task; check_ans;
	give_id_245; give_act_reap; latency_task; check_ans;
	give_id_246; give_act_reap; latency_task; check_ans;
	give_id_247; give_act_reap; latency_task; check_ans;
	give_id_248; give_act_reap; latency_task; check_ans;
	give_id_249; give_act_reap; latency_task; check_ans;
	give_id_250; give_act_reap; latency_task; check_ans;
	give_id_251; give_act_reap; latency_task; check_ans;
	give_id_252; give_act_reap; latency_task; check_ans;
	give_id_253; give_act_reap; latency_task; check_ans;
	give_id_254; give_act_reap; latency_task; check_ans;


    // for(user_num=0; user_num < user_num ; user_num = user_num +1)begin
		// input_task;
		// wait_out_valid;
		// check_ans;
		// repeat(3) @(negedge clk);
    // end
	// input_task;
	// #(2000);
	congratulations;
	// $finish;
end

// initial begin
	// #(1000);
	// $finish;
	// congratulations;
// end

// initial begin
	// forever@(posedge clk)begin
		// if(inf.out_valid)begin
		    // @(negedge clk);
			// if((inf.complete    !== golden_complete) ||
			   // (inf.err_msg     !== golden_err_msg ) ||
			   // (inf.out_info    !== golden_out_info) ||
			   // (inf.out_deposit !== golden_out_deposit) ) begin
				// #(100)
				// $finish;
			// end
            // else begin

				// $display("\033[0;38;5;111mPASS USER \033[4m NO.%3d \033[m \033[0;38;5;219mACT NO. %d\033[m latency: %3d", user_cnt, act_cnt, wait_val_time);
            // end			
		// end
	// end
// end

//================================================================
// task definition
//================================================================
task reset_signal_task; begin 
    #(0.5);  inf.rst_n <= 0;
    $readmemh(DRAM_p_r, golden_DRAM);	
	inf.D           = 0;
	inf.id_valid    = 0;
	inf.cat_valid   = 0;
	inf.amnt_valid  = 0;
	inf.act_valid   = 0;
	#(5);
	if((inf.out_valid   !== 'b0)||
	   (inf.complete    !== 'b0)||
	   (inf.err_msg     !== 'b0)||
	   (inf.out_info    !== 'b0)||
	   (inf.out_deposit !== 'b0)) begin
		// $display("************************************************************");
		// $display("*                             FAIL                         *");
		// $display("*   Output signal should be 0 after initial RESET at %t    *",$time);
		// $display("************************************************************");
		// $finish;
	end
    #(5);
	inf.rst_n <=1;
end endtask

task latency_task; begin 
    lat=-1;
    while(inf.out_valid!==1) begin
		lat=lat+1;
		if(lat==1200)begin
			// if(lat==50)begin
				// $display ("*********************************************************");
				// $display ("*                     SPEC 6 FAIL!                      *");
				// $display ("*       The execution latency are over 300 cycles.      *");
				// $display ("*********************************************************");
				// $display("  SPEC 6 FAIL!  ");
			// end
			// repeat(2)@(negedge clk);
			// $finish;
		end
		@(negedge clk);
    end
	// @(negedge clk);
	total_latency = total_latency + lat;
end endtask

task input_task; begin
    // D,
	// id_valid,
	// passwd_valid,
	// amnt_valid,
	// act_valid,
	// C_out_valid,
	// C_data_r
	
	// user_log_in;
	// r_act.randomize();
	// case(r_act.ran_act)
		// 3'd2:
		// 3'd3:
		// 3'd5:
		// 3'd6:
		// 3'd7:
	// endcase
	
	//transfer_money;
	// make_a_deposit;
	//check_balance;
    //change_user_password;
	
    // user_log_out;
	// user_log_in;
end
endtask
task check_ans; begin
	// $display("golden_id = %d",golden_id);
	// 0~255 -> 65536~66559(66560)
	// $display("land id = %d",golden_DRAM[golden_id+65536]);
	// $display("land crop = %d",golden_DRAM[golden_id+65536+1][3:0]);
	// $display("land status = %d",golden_DRAM[golden_id+65536+1][7:4]);
	// $display("land water = %d",golden_DRAM[golden_id+65536+2]);
	// $display("land water = %d",golden_DRAM[golden_id+65536+3]);
	// golden_land_info.land_id     = golden_DRAM[golden_id+65536];
	// golden_land_info.land_status = golden_DRAM[golden_id+65536+1];
	// golden_land_info.water_amnt  = {golden_DRAM[golden_id+65536+2],golden_DRAM[golden_id+65536+3]};
	// $display("land id = %d",golden_land_info.land_id);
	// $display("land crop = %d",golden_land_info.land_status);
	// $display("land water = %d",golden_land_info.water_amnt);
	golden_land_id     = golden_DRAM[golden_id*4+65536];
	golden_land_crop   = golden_DRAM[golden_id*4+65536+1][3:0];
	golden_land_status = golden_DRAM[golden_id*4+65536+1][7:4];
	golden_land_water  = {golden_DRAM[golden_id*4+65536+2],golden_DRAM[golden_id*4+65536+3]};
	// $display("golden_land_water = %d",golden_land_water);
	
	if ((golden_act == Seed) && ((golden_land_status == Zer_sta) || (golden_land_status == Fst_sta) || (golden_land_status == Snd_sta))) begin
		golden_complete = 0;
		golden_err_msg = Not_Empty;
	end
	else if ((golden_act == Water) && (golden_land_status == No_sta)) begin
		golden_complete = 0;
		golden_err_msg = Is_Empty;
	end
	else if ((golden_act == Water) && (golden_land_status == Snd_sta)) begin
		golden_complete = 0;
		golden_err_msg = Has_Grown;
	end
	else if ((golden_act == Reap) && (golden_land_status == No_sta)) begin
		golden_complete = 0;
		golden_err_msg = Is_Empty;
	end
	else if ((golden_act == Reap) && (golden_land_status == Zer_sta)) begin
		golden_complete = 0;
		golden_err_msg = Not_Grown;
	end
	else if ((golden_act == Steal) && (golden_land_status == No_sta)) begin
		golden_complete = 0;
		golden_err_msg = Is_Empty;
	end
	else if ((golden_act == Steal) && (golden_land_status == Zer_sta)) begin
		golden_complete = 0;
		golden_err_msg = Not_Grown;
	end
	else begin
		golden_complete = 1;
		golden_err_msg = No_Err;
	end
		
	if (golden_complete == 1) begin
		if (golden_act == Seed) begin
			if ((golden_land_status == No_sta) || (golden_land_status == 0)) begin
				golden_land_crop   = golden_crop;
				// golden_land_status = Zer_sta;
				golden_land_water  = golden_land_water + golden_water;
				case (golden_land_crop)
					Potato: begin
						golden_deposit = golden_deposit - 'd5;
						if (golden_land_water >= 16'h0080)
							golden_land_status = Snd_sta;
						else if (golden_land_water >= 16'h0010)
							golden_land_status = Fst_sta;
						else
							golden_land_status = Zer_sta;
					end
					Corn: begin
						golden_deposit = golden_deposit - 'd10;
						if (golden_land_water >= 16'h0200)
							golden_land_status = Snd_sta;
						else if (golden_land_water >= 16'h0040)
							golden_land_status = Fst_sta;
						else
							golden_land_status = Zer_sta;
					end
					Tomato: begin
						golden_deposit = golden_deposit - 'd15;
						if (golden_land_water >= 16'h0800)
							golden_land_status = Snd_sta;
						else if (golden_land_water >= 16'h0100)
							golden_land_status = Fst_sta;
						else
							golden_land_status = Zer_sta;
					end
					Wheat: begin
						golden_deposit = golden_deposit - 'd20;
						if (golden_land_water >= 16'h2000)
							golden_land_status = Snd_sta;
						else if (golden_land_water >= 16'h0400)
							golden_land_status = Fst_sta;
						else
							golden_land_status = Zer_sta;
					end
				endcase
			end
			golden_out_info = {golden_land_id,golden_land_status,golden_land_crop,golden_land_water};
			golden_out_deposit = 0;
		end
		else if (golden_act == Water) begin
			if ((golden_land_status == Zer_sta) || (golden_land_status == Fst_sta))
				golden_land_water  = golden_land_water + golden_water;
			case (golden_land_crop)
				Potato: begin
					if (golden_land_water >= 16'h0080)
						golden_land_status = Snd_sta;
					else if (golden_land_water >= 16'h0010)
						golden_land_status = Fst_sta;
					else
						golden_land_status = Zer_sta;
				end
				Corn: begin
					if (golden_land_water >= 16'h0200)
						golden_land_status = Snd_sta;
					else if (golden_land_water >= 16'h0040)
						golden_land_status = Fst_sta;
					else
						golden_land_status = Zer_sta;
				end
				Tomato: begin
					if (golden_land_water >= 16'h0800)
						golden_land_status = Snd_sta;
					else if (golden_land_water >= 16'h0100)
						golden_land_status = Fst_sta;
					else
						golden_land_status = Zer_sta;
				end
				Wheat: begin
					if (golden_land_water >= 16'h2000)
						golden_land_status = Snd_sta;
					else if (golden_land_water >= 16'h0400)
						golden_land_status = Fst_sta;
					else
						golden_land_status = Zer_sta;
				end
			endcase
			golden_out_info = {golden_land_id,golden_land_status,golden_land_crop,golden_land_water};
			golden_out_deposit = 0;
		end
		else if (golden_act == Reap) begin
			// if ((golden_land_status == Fst_sta) || (golden_land_status == Snd_sta)) begin
				// golden_deposit = golden_deposit - 'd5;
				// if (golden_land_status == Fst_sta) begin
					// case (golden_land_crop)
						// Potato: deposit = deposit + 'd10;
						// Corn  : deposit = deposit + 'd20;
						// Tomato: deposit = deposit + 'd30;
						// Wheat : deposit = deposit + 'd40;
					// endcase
				// end
				// else if (golden_land_status == Snd_sta) begin
					// case (golden_land_crop)
						// Potato: deposit = deposit + 'd25;
						// Corn  : deposit = deposit + 'd50;
						// Tomato: deposit = deposit + 'd75;
						// Wheat : deposit = deposit + 'd100;
					// endcase
				// end
				// golden_land_status = No_sta;
				// golden_land_water  = 0;
			// end
			golden_out_info = {golden_land_id,golden_land_status,golden_land_crop,golden_land_water};
			golden_out_deposit = 0;
		end
		else if (golden_act == Steal) begin
			// if ((golden_land_status == Fst_sta) || (golden_land_status == Snd_sta)) begin
				// golden_land_status = No_sta;
				// golden_land_water  = 0;
			// end
			golden_out_info = {golden_land_id,golden_land_status,golden_land_crop,golden_land_water};
			golden_out_deposit = 0;
		end
		else if (golden_act == Check_dep) begin
			golden_out_info = 0;
			golden_out_deposit = golden_deposit;
		end
	end
	else begin // golden_complete == 0
		golden_out_info = 0;
		golden_out_deposit = 0;
	end
	// golden_out_info = {golden_land_id,golden_land_status,golden_land_crop,golden_land_water};
	// golden_out_deposit = 0;
	if ((golden_complete    !== inf.complete)    ||
	    (golden_err_msg     !== inf.err_msg)     ||
	    (golden_out_info    !== inf.out_info)    ||
	    (golden_out_deposit !== inf.out_deposit)) begin
		$display("*********************************************************************");
		$display("*                             FAIL!                                 *");		
		$display("*    golden_complete    : %8d,  Your complete    : %8d    *",golden_complete   ,inf.complete);
		$display("*    golden_err_msg     : %8d,  Your err_msg     : %8d    *",golden_err_msg    ,inf.err_msg);
		$display("*    golden_out_info    : %8h,  Your out_info    : %8h    *",golden_out_info   ,inf.out_info);
		$display("*    golden_out_deposit : %8h,  Your out_deposit : %8h    *",golden_out_deposit,inf.out_deposit);
		$display("*********************************************************************");
		repeat(2) @(negedge clk);
		$finish;
	end
	
	if (golden_complete == 1) begin
		if (golden_act == Reap) begin
			if ((golden_land_status == Fst_sta) || (golden_land_status == Snd_sta)) begin
				// golden_deposit = golden_deposit - 'd5;
				if (golden_land_status == Fst_sta) begin
					case (golden_land_crop)
						Potato: golden_deposit = golden_deposit + 'd10;
						Corn  : golden_deposit = golden_deposit + 'd20;
						Tomato: golden_deposit = golden_deposit + 'd30;
						Wheat : golden_deposit = golden_deposit + 'd40;
					endcase
				end
				else if (golden_land_status == Snd_sta) begin
					case (golden_land_crop)
						Potato: golden_deposit = golden_deposit + 'd25;
						Corn  : golden_deposit = golden_deposit + 'd50;
						Tomato: golden_deposit = golden_deposit + 'd75;
						Wheat : golden_deposit = golden_deposit + 'd100;
					endcase
				end
				golden_land_status = No_sta;
				golden_land_water  = 0;
			end
		end
		else if (golden_act == Steal) begin
			if ((golden_land_status == Fst_sta) || (golden_land_status == Snd_sta)) begin
				golden_land_status = No_sta;
				golden_land_water  = 0;
			end
		end
	end
	
	golden_DRAM[golden_id*4+65536] = golden_land_id;
	golden_DRAM[golden_id*4+65536+1][3:0] = golden_land_crop;
	golden_DRAM[golden_id*4+65536+1][7:4] = golden_land_status;
	golden_DRAM[golden_id*4+65536+2] = golden_land_water[15:8];
	golden_DRAM[golden_id*4+65536+3] = golden_land_water[ 7:0];
	
	@(negedge clk);
end
endtask

task give_id; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.randomize();
	golden_id = r_id.ran_id;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_0; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(0);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
	// $display("%d",golden_id);
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_1; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(1);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_2; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(2);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_3; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(3);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_4; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(4);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_5; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(5);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_6; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(6);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_7; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(7);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_8; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(8);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_9; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(9);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_10; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(10);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_11; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(11);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_12; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(12);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_13; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(13);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_14; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(14);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_15; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(15);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_16; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(16);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_17; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(17);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_18; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(18);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_19; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(19);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_20; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(20);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_21; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(21);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_22; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(22);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_23; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(23);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_24; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(24);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_25; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(25);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_26; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(26);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_27; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(27);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_28; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(28);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_29; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(29);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_30; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(30);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_31; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(31);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_32; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(32);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_33; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(33);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_34; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(34);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_35; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(35);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_36; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(36);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_37; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(37);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_38; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(38);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_39; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(39);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_40; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(40);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_41; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(41);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_42; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(42);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_43; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(43);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_44; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(44);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_45; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(45);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_46; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(46);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_47; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(47);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_48; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(48);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_49; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(49);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_50; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(50);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_51; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(51);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_52; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(52);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_53; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(53);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_54; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(54);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_55; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(55);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_56; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(56);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_57; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(57);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_58; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(58);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_59; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(59);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_60; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(60);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_61; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(61);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_62; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(62);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_63; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(63);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_64; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(64);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_65; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(65);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_66; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(66);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_67; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(67);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_68; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(68);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_69; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(69);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_70; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(70);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_71; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(71);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_72; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(72);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_73; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(73);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_74; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(74);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_75; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(75);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_76; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(76);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_77; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(77);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_78; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(78);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_79; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(79);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_80; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(80);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_81; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(81);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_82; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(82);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_83; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(83);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_84; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(84);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_85; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(85);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_86; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(86);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_87; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(87);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_88; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(88);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_89; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(89);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_90; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(90);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_91; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(91);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_92; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(92);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_93; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(93);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_94; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(94);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_95; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(95);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_96; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(96);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_97; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(97);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_98; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(98);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_99; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(99);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_100; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(100);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_101; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(101);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_102; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(102);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_103; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(103);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_104; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(104);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_105; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(105);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_106; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(106);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_107; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(107);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_108; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(108);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_109; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(109);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_110; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(110);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_111; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(111);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_112; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(112);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_113; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(113);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_114; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(114);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_115; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(115);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_116; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(116);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_117; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(117);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_118; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(118);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_119; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(119);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_120; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(120);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_121; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(121);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_122; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(122);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_123; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(123);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_124; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(124);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_125; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(125);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_126; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(126);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_127; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(127);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_128; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(128);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_129; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(129);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_130; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(130);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_131; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(131);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_132; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(132);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_133; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(133);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_134; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(134);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_135; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(135);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_136; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(136);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_137; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(137);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_138; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(138);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_139; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(139);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_140; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(140);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_141; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(141);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_142; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(142);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_143; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(143);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_144; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(144);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_145; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(145);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_146; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(146);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_147; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(147);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_148; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(148);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_149; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(149);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_150; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(150);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_151; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(151);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_152; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(152);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_153; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(153);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_154; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(154);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_155; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(155);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_156; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(156);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_157; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(157);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_158; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(158);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_159; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(159);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_160; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(160);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_161; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(161);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_162; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(162);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_163; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(163);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_164; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(164);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_165; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(165);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_166; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(166);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_167; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(167);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_168; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(168);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_169; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(169);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_170; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(170);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_171; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(171);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_172; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(172);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_173; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(173);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_174; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(174);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_175; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(175);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_176; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(176);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_177; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(177);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_178; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(178);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_179; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(179);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_180; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(180);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_181; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(181);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_182; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(182);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_183; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(183);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_184; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(184);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_185; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(185);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_186; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(186);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_187; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(187);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_188; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(188);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_189; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(189);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_190; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(190);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_191; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(191);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_192; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(192);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_193; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(193);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_194; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(194);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_195; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(195);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_196; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(196);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_197; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(197);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_198; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(198);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_199; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(199);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_200; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(200);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_201; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(201);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_202; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(202);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_203; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(203);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_204; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(204);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_205; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(205);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_206; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(206);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_207; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(207);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_208; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(208);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_209; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(209);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_210; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(210);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_211; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(211);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_212; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(212);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_213; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(213);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_214; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(214);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_215; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(215);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_216; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(216);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_217; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(217);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_218; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(218);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_219; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(219);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_220; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(220);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_221; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(221);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_222; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(222);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_223; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(223);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_224; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(224);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_225; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(225);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_226; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(226);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_227; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(227);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_228; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(228);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_229; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(229);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_230; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(230);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_231; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(231);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_232; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(232);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_233; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(233);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_234; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(234);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_235; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(235);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_236; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(236);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_237; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(237);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_238; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(238);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_239; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(239);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_240; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(240);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_241; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(241);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_242; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(242);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_243; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(243);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_244; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(244);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_245; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(245);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_246; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(246);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_247; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(247);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_248; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(248);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_249; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(249);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_250; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(250);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_251; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(251);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_252; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(252);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_253; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(253);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_254; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(254);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask

task give_id_255; begin
	repeat(1) @(negedge clk);
	inf.id_valid = 'b1;
	r_id.set(255);
	golden_id = r_id.out;
	inf.D     = {8'b0, golden_id};
    repeat(1) @(negedge clk);
	inf.id_valid = 'b0;
	inf.D        = 'dx;
end
endtask


task give_act; begin
	repeat(1) @(negedge clk);
	inf.act_valid = 'b1;
	r_act.randomize();
	golden_act = r_act.ran_act;
	inf.D     = {12'b0, golden_act};
    repeat(1) @(negedge clk);
	inf.act_valid = 'b0;
	inf.D         = 'dx;
end
endtask

task give_act_seed; begin
	// act_valid
	repeat(1) @(negedge clk);
	inf.act_valid = 'b1;
	golden_act = Seed;
	inf.D     = {12'b0, golden_act};
    repeat(1) @(negedge clk);
	inf.act_valid = 'b0;
	inf.D         = 'dx;
	// cat_valid
	repeat(1) @(negedge clk);
	inf.cat_valid = 'b1;
	r_crop.randomize();
	golden_crop = r_crop.ran_crop;
	inf.D       = {12'b0, golden_crop};
    repeat(1) @(negedge clk);
	inf.cat_valid = 'b0;
	inf.D         = 'dx;
	// amnt_valid
	repeat(1) @(negedge clk);
	inf.amnt_valid = 'b1;
	r_water.randomize();
	golden_water = r_water.ran_water;
	inf.D       = {golden_water};
    repeat(1) @(negedge clk);
	inf.amnt_valid = 'b0;
	inf.D          = 'dx;
end
endtask

task give_act_seed_actual_0; begin
	// act_valid
	repeat(1) @(negedge clk);
	inf.act_valid = 'b1;
	golden_act = Seed;
	inf.D     = {12'b0, golden_act};
    repeat(1) @(negedge clk);
	inf.act_valid = 'b0;
	inf.D         = 'dx;
	// cat_valid
	repeat(1) @(negedge clk);
	inf.cat_valid = 'b1;
	r_crop.randomize();
	golden_crop = r_crop.ran_crop;
	inf.D       = {12'b0, golden_crop};
    repeat(1) @(negedge clk);
	inf.cat_valid = 'b0;
	inf.D         = 'dx;
	// amnt_valid
	repeat(1) @(negedge clk);
	inf.amnt_valid = 'b1;
	golden_water = 16'd0;
	inf.D       = {golden_water};
    repeat(1) @(negedge clk);
	inf.amnt_valid = 'b0;
	inf.D          = 'dx;
end
endtask

task give_act_seed_water_1; begin
	// act_valid
	repeat(1) @(negedge clk);
	inf.act_valid = 'b1;
	golden_act = Seed;
	inf.D     = {12'b0, golden_act};
    repeat(1) @(negedge clk);
	inf.act_valid = 'b0;
	inf.D         = 'dx;
	// cat_valid
	repeat(1) @(negedge clk);
	inf.cat_valid = 'b1;
	r_crop.randomize();
	golden_crop = r_crop.ran_crop;
	inf.D       = {12'b0, golden_crop};
    repeat(1) @(negedge clk);
	inf.cat_valid = 'b0;
	inf.D         = 'dx;
	// amnt_valid
	repeat(1) @(negedge clk);
	inf.amnt_valid = 'b1;
	r_water.randomize();
	golden_water = r_water.ran_water_1;
	inf.D       = {golden_water};
    repeat(1) @(negedge clk);
	inf.amnt_valid = 'b0;
	inf.D          = 'dx;
end
endtask

task give_crop; begin
	repeat(1) @(negedge clk);
	inf.cat_valid = 'b1;
	r_crop.randomize();
	golden_crop = r_crop.ran_crop;
	inf.D       = {12'b0, golden_crop};
    repeat(1) @(negedge clk);
	inf.cat_valid = 'b0;
	inf.D         = 'dx;
end
endtask

task give_water; begin
	repeat(1) @(negedge clk);
	inf.act_valid = 'b1;
	golden_act = Water;
	inf.D      = {12'b0, golden_act};
	repeat(1) @(negedge clk);
	inf.act_valid = 'b0;
	inf.D         = 'dx;
	repeat(1) @(negedge clk);
	inf.amnt_valid = 'b1;
	r_water.randomize();
	golden_water = r_water.ran_water;
	inf.D       = {golden_water};
    repeat(1) @(negedge clk);
	inf.amnt_valid = 'b0;
	inf.D          = 'dx;
end
endtask

task give_water_0; begin
	repeat(1) @(negedge clk);
	inf.act_valid = 'b1;
	golden_act = Water;
	inf.D      = {12'b0, golden_act};
	repeat(1) @(negedge clk);
	inf.act_valid = 'b0;
	inf.D         = 'dx;
	repeat(1) @(negedge clk);
	inf.amnt_valid = 'b1;
	r_water.randomize();
	golden_water = r_water.ran_water_0;
	// $display("%d",golden_water);
	inf.D       = {golden_water};
    repeat(1) @(negedge clk);
	inf.amnt_valid = 'b0;
	inf.D          = 'dx;
end
endtask

task give_water_1; begin
	repeat(1) @(negedge clk);
	inf.act_valid = 'b1;
	golden_act = Water;
	inf.D      = {12'b0, golden_act};
	repeat(1) @(negedge clk);
	inf.act_valid = 'b0;
	inf.D         = 'dx;
	repeat(1) @(negedge clk);
	inf.amnt_valid = 'b1;
	r_water.randomize();
	golden_water = r_water.ran_water_1;
	inf.D       = {golden_water};
    repeat(1) @(negedge clk);
	inf.amnt_valid = 'b0;
	inf.D          = 'dx;
end
endtask
task give_water_2; begin
	repeat(1) @(negedge clk);
	inf.act_valid = 'b1;
	golden_act = Water;
	inf.D      = {12'b0, golden_act};
	repeat(1) @(negedge clk);
	inf.act_valid = 'b0;
	inf.D         = 'dx;
	repeat(1) @(negedge clk);
	inf.amnt_valid = 'b1;
	r_water.randomize();
	golden_water = r_water.ran_water_2;
	inf.D       = {golden_water};
    repeat(1) @(negedge clk);
	inf.amnt_valid = 'b0;
	inf.D          = 'dx;
end
endtask

task give_water_3; begin
	repeat(1) @(negedge clk);
	inf.act_valid = 'b1;
	golden_act = Water;
	inf.D      = {12'b0, golden_act};
	repeat(1) @(negedge clk);
	inf.act_valid = 'b0;
	inf.D         = 'dx;
	repeat(1) @(negedge clk);
	inf.amnt_valid = 'b1;
	r_water.randomize();
	golden_water = r_water.ran_water_3;
	inf.D       = {golden_water};
    repeat(1) @(negedge clk);
	inf.amnt_valid = 'b0;
	inf.D          = 'dx;
end
endtask

task give_water_4; begin
	repeat(1) @(negedge clk);
	inf.act_valid = 'b1;
	golden_act = Water;
	inf.D      = {12'b0, golden_act};
	repeat(1) @(negedge clk);
	inf.act_valid = 'b0;
	inf.D         = 'dx;
	repeat(1) @(negedge clk);
	inf.amnt_valid = 'b1;
	r_water.randomize();
	golden_water = r_water.ran_water_4;
	inf.D       = {golden_water};
    repeat(1) @(negedge clk);
	inf.amnt_valid = 'b0;
	inf.D          = 'dx;
end
endtask

task give_water_5; begin
	repeat(1) @(negedge clk);
	inf.act_valid = 'b1;
	golden_act = Water;
	inf.D      = {12'b0, golden_act};
	repeat(1) @(negedge clk);
	inf.act_valid = 'b0;
	inf.D         = 'dx;
	repeat(1) @(negedge clk);
	inf.amnt_valid = 'b1;
	r_water.randomize();
	golden_water = r_water.ran_water_5;
	inf.D       = {golden_water};
    repeat(1) @(negedge clk);
	inf.amnt_valid = 'b0;
	inf.D          = 'dx;
end
endtask

task give_water_actual_0; begin
	repeat(1) @(negedge clk);
	inf.act_valid = 'b1;
	golden_act = Water;
	inf.D      = {12'b0, golden_act};
	repeat(1) @(negedge clk);
	inf.act_valid = 'b0;
	inf.D         = 'dx;
	repeat(1) @(negedge clk);
	inf.amnt_valid = 'b1;
	golden_water = 16'd0;
	inf.D       = {golden_water};
    repeat(1) @(negedge clk);
	inf.amnt_valid = 'b0;
	inf.D          = 'dx;
end
endtask

task give_act_reap; begin
	repeat(1) @(negedge clk);
	inf.act_valid = 'b1;
	golden_act = Reap;
	inf.D     = {12'b0, golden_act};
    repeat(1) @(negedge clk);
	inf.act_valid = 'b0;
	inf.D         = 'dx;
end
endtask

task give_act_steal; begin
	repeat(1) @(negedge clk);
	inf.act_valid = 'b1;
	golden_act = Steal;
	inf.D     = {12'b0, golden_act};
    repeat(1) @(negedge clk);
	inf.act_valid = 'b0;
	inf.D         = 'dx;
end
endtask

task give_check_deposit; begin
	repeat(1) @(negedge clk);
	inf.act_valid = 'b1;
	golden_act = Check_dep;
	inf.D         = {12'b0, golden_act};
    repeat(1) @(negedge clk);
	inf.act_valid = 'b0;
	inf.D         = 'dx;
end
endtask

task congratulations; begin
    $display("********************************************************************");
    $display("                        \033[0;38;5;219mCongratulations!\033[m      ");
    $display("                 \033[0;38;5;219mYou have passed all patterns!\033[m");
    $display("                 \033[0;38;5;219mTotal time: %d \033[m",$time);
    $display("********************************************************************");
    // image_.success;
	repeat(2) @(negedge clk);
    $finish;
end
endtask

endprogram


