module CHIP(
    clk,
    rst_n,
    in_valid,
    in_data,
    size,
    action,
    out_valid,
    out_data
);

input [31:0] in_data;
input [1:0] size;
input [2:0] action;
input clk, rst_n, in_valid;

output [31:0] out_data;
output out_valid;

wire C_clk, C_in_valid, C_rst_n;
wire [31:0] C_in_data,C_out_data;
wire [1:0] C_size;
wire [2:0] C_action;
wire BUF_CLK;
// TA has already defined for you
// MC module
MC MC (
    .clk(BUF_CLK),
    .rst_n(C_rst_n),
    .in_valid(C_in_valid),
    .in_data(C_in_data),
    .size(C_size),
    .action(C_action),
    .out_valid(C_out_valid),
    .out_data(C_out_data)
);

CLKBUFX20 buf0(.A(C_clk),.Y(BUF_CLK));

P8C I_CLK      ( .Y(C_clk),         .P(clk),         .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b0), .CSEN(1'b1) );
P8C I_RESET    ( .Y(C_rst_n),       .P(rst_n),       .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_VALID    ( .Y(C_in_valid),    .P(in_valid),    .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_SIZE_0   ( .Y(C_size[0]),     .P(size[0]),     .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_SIZE_1   ( .Y(C_size[1]),     .P(size[1]),     .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_ACTION_0 ( .Y(C_action[0]),   .P(action[0]),   .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_ACTION_1 ( .Y(C_action[1]),   .P(action[1]),   .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_ACTION_2 ( .Y(C_action[2]),   .P(action[2]),   .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_0     ( .Y(C_in_data[0 ]), .P(in_data[0 ]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_1     ( .Y(C_in_data[1 ]), .P(in_data[1 ]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_2     ( .Y(C_in_data[2 ]), .P(in_data[2 ]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_3     ( .Y(C_in_data[3 ]), .P(in_data[3 ]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_4     ( .Y(C_in_data[4 ]), .P(in_data[4 ]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_5     ( .Y(C_in_data[5 ]), .P(in_data[5 ]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_6     ( .Y(C_in_data[6 ]), .P(in_data[6 ]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_7     ( .Y(C_in_data[7 ]), .P(in_data[7 ]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_8     ( .Y(C_in_data[8 ]), .P(in_data[8 ]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_9     ( .Y(C_in_data[9 ]), .P(in_data[9 ]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_10    ( .Y(C_in_data[10]), .P(in_data[10]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_11    ( .Y(C_in_data[11]), .P(in_data[11]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_12    ( .Y(C_in_data[12]), .P(in_data[12]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_13    ( .Y(C_in_data[13]), .P(in_data[13]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_14    ( .Y(C_in_data[14]), .P(in_data[14]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_15    ( .Y(C_in_data[15]), .P(in_data[15]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_16    ( .Y(C_in_data[16]), .P(in_data[16]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_17    ( .Y(C_in_data[17]), .P(in_data[17]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_18    ( .Y(C_in_data[18]), .P(in_data[18]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_19    ( .Y(C_in_data[19]), .P(in_data[19]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_20    ( .Y(C_in_data[20]), .P(in_data[20]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_21    ( .Y(C_in_data[21]), .P(in_data[21]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_22    ( .Y(C_in_data[22]), .P(in_data[22]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_23    ( .Y(C_in_data[23]), .P(in_data[23]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_24    ( .Y(C_in_data[24]), .P(in_data[24]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_25    ( .Y(C_in_data[25]), .P(in_data[25]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_26    ( .Y(C_in_data[26]), .P(in_data[26]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_27    ( .Y(C_in_data[27]), .P(in_data[27]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_28    ( .Y(C_in_data[28]), .P(in_data[28]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_29    ( .Y(C_in_data[29]), .P(in_data[29]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_30    ( .Y(C_in_data[30]), .P(in_data[30]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_31    ( .Y(C_in_data[31]), .P(in_data[31]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );

P8C O_VALID    ( .A(C_out_valid), 	 .P(out_valid),    .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_0    ( .A(C_out_data[0 ]), .P(out_data[0 ]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_1    ( .A(C_out_data[1 ]), .P(out_data[1 ]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_2    ( .A(C_out_data[2 ]), .P(out_data[2 ]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_3    ( .A(C_out_data[3 ]), .P(out_data[3 ]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_4    ( .A(C_out_data[4 ]), .P(out_data[4 ]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_5    ( .A(C_out_data[5 ]), .P(out_data[5 ]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_6    ( .A(C_out_data[6 ]), .P(out_data[6 ]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_7    ( .A(C_out_data[7 ]), .P(out_data[7 ]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_8    ( .A(C_out_data[8 ]), .P(out_data[8 ]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_9    ( .A(C_out_data[9 ]), .P(out_data[9 ]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_10   ( .A(C_out_data[10]), .P(out_data[10]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_11   ( .A(C_out_data[11]), .P(out_data[11]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_12   ( .A(C_out_data[12]), .P(out_data[12]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_13   ( .A(C_out_data[13]), .P(out_data[13]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_14   ( .A(C_out_data[14]), .P(out_data[14]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_15   ( .A(C_out_data[15]), .P(out_data[15]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_16   ( .A(C_out_data[16]), .P(out_data[16]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_17   ( .A(C_out_data[17]), .P(out_data[17]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_18   ( .A(C_out_data[18]), .P(out_data[18]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_19   ( .A(C_out_data[19]), .P(out_data[19]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_20   ( .A(C_out_data[20]), .P(out_data[20]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_21   ( .A(C_out_data[21]), .P(out_data[21]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_22   ( .A(C_out_data[22]), .P(out_data[22]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_23   ( .A(C_out_data[23]), .P(out_data[23]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_24   ( .A(C_out_data[24]), .P(out_data[24]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_25   ( .A(C_out_data[25]), .P(out_data[25]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_26   ( .A(C_out_data[26]), .P(out_data[26]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_27   ( .A(C_out_data[27]), .P(out_data[27]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_28   ( .A(C_out_data[28]), .P(out_data[28]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_29   ( .A(C_out_data[29]), .P(out_data[29]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_30   ( .A(C_out_data[30]), .P(out_data[30]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_31   ( .A(C_out_data[31]), .P(out_data[31]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));

// I/O power 3.3V pads x? (DVDD + DGND) 40 output 33 input
PVDDR VDDP0  (); PVSSR GNDP0  ();
PVDDR VDDP1  (); PVSSR GNDP1  ();
PVDDR VDDP2  (); PVSSR GNDP2  ();
PVDDR VDDP3  (); PVSSR GNDP3  ();
PVDDR VDDP4  (); PVSSR GNDP4  ();
PVDDR VDDP5  (); PVSSR GNDP5  ();
PVDDR VDDP6  (); PVSSR GNDP6  ();
PVDDR VDDP7  (); PVSSR GNDP7  ();
// PVDDR VDDP8  (); PVSSR GNDP8  ();
// PVDDR VDDP9  (); PVSSR GNDP9  ();
// PVDDR VDDP10 (); PVSSR GNDP10 ();
// PVDDR VDDP11 (); PVSSR GNDP11 ();
// PVDDR VDDP12 (); PVSSR GNDP12 ();
// PVDDR VDDP13 (); PVSSR GNDP13 ();


// Core poweri 1.8V pads x? (VDD + GND) 40 output 33 input
PVDDC VDDC0  (); PVSSC GNDC0  ();
PVDDC VDDC1  (); PVSSC GNDC1  ();
PVDDC VDDC2  (); PVSSC GNDC2  ();
PVDDC VDDC3  (); PVSSC GNDC3  ();
PVDDC VDDC4  (); PVSSC GNDC4  ();
PVDDC VDDC5  (); PVSSC GNDC5  ();
PVDDC VDDC6  (); PVSSC GNDC6  ();
PVDDC VDDC7  (); PVSSC GNDC7  ();
// PVDDC VDDC8  (); PVSSC GNDC8  ();
// PVDDC VDDC9  (); PVSSC GNDC9  ();
// PVDDC VDDC10 (); PVSSC GNDC10 ();
// PVDDC VDDC11 (); PVSSC GNDC11 ();
// PVDDC VDDC12 (); PVSSC GNDC12 ();
// PVDDC VDDC13 (); PVSSC GNDC13 ();

endmodule
